* SPICE NETLIST
***************************************

.SUBCKT pvar18_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar33_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rnwaa_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rnwsti_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rpdif_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rndif_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rppo_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rppo_3t_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rnpo_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rnpo_3t_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rpdifsab_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rndifsab_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rpposab_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rpposab_3t_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rnposab_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rnposab_3t_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT rhrpo_ckt PLUS MINUS
.ENDS
***************************************
.SUBCKT rhrpo_3t_ckt PLUS MINUS SUB
.ENDS
***************************************
.SUBCKT n18_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw18_ckt_rf DRN GATE SRC BULK T
.ENDS
***************************************
.SUBCKT p18_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT n33_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT dnw33_ckt_rf DRN GATE SRC BULK T
.ENDS
***************************************
.SUBCKT p33_ckt_rf DRN GATE SRC BULK
.ENDS
***************************************
.SUBCKT pvar18w10l1_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18w10ld5_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18w5l1_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar18w5ld5_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar33w10l1_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvar33w10ld5_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvardio18_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT pvardio33_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rndifsab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rpdifsab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rnposab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rpposab_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT rhrpo_ckt_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mim1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT ind_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT diff_ind_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT diff_ind_3t_rf PLUS MINUS B
.ENDS
***************************************
