*****************************************************************************
* CDL NETLIST:
* CELL NAME: ALL_CELL
* NETLISTED ON: AUG 20 14:51:26 2004
*****************************************************************************


*****************************************************************************
* GLOBAL NET DECLARATIONS
*****************************************************************************
*.GLOBAL VDD GND


*****************************************************************************
* PIN CONTROL STATEMENT
*****************************************************************************
*.PIN VDD GND


*****************************************************************************
* BIPOLAR DECLARATIONS
*****************************************************************************


*.BIPOLAR
*.RESI = 1.000000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.SCALE METER
*.LDD

*****************************************************************************
* PARAMETER STATEMENT
*****************************************************************************
.PARAM


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TG1G                                                                 *
* LAST TIME SAVED: SEP 10 14:41:27 2001                                       *
*******************************************************************************
.SUBCKT TG1G D Q CK CKB NL=0.18U NW=0.24U PL=0.18U PW=0.24U
*.NOPIN VDD GND
MP0 Q CKB D VDD P18 W=PW L=PL
MN0 D CK Q GND N18 W=NW L=NL
.ENDS TG1G


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IVG                                                                  *
* LAST TIME SAVED: SEP 10 14:37:09 2001                                       *
*******************************************************************************
.SUBCKT IVG Z A PL=0.18U PW=0.24U NL=0.18U NW=0.24U
MN0 Z A GND GND N18 W=NW L=NL
MP0 VDD A Z VDD P18 W=PW L=PL
.ENDS IVG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR3HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:45:44 2002                                       *
*******************************************************************************
.SUBCKT XOR3HD4X Z A B C
XI8 NET13 NET21 NET17 B TG1G NW=2U PW=2U
XI9 NET15 NET21 B NET17 TG1G NW=2U PW=2U
XI5 NET13 NET29 B NET17 TG1G NW=2U PW=2U
XI3 NET15 NET29 NET17 B TG1G NW=2U PW=2U
XI4 NET21 NET6 NET35 C TG1G NW=2U PW=2U
XI2 NET29 NET6 C NET35 TG1G NW=2U PW=2U
XI10 NET35 C IVG PW=0.9U NW=0.6U
XI7 NET13 A IVG PW=3.44U NW=2.4U
XI6 NET15 NET13 IVG PW=3.44U NW=2.4U
XI0 NET17 B IVG PW=1.68U NW=1.18U
XI1 Z NET6 IVG PW=4.8U NW=3.2U
.ENDS XOR3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR3HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:45:40 2002                                       *
*******************************************************************************
.SUBCKT XOR3HD2X Z A B C
XI8 NET13 NET21 NET17 B TG1G NW=1.18U PW=1.18U
XI9 NET15 NET21 B NET17 TG1G NW=1.18U PW=1.18U
XI5 NET13 NET29 B NET17 TG1G NW=1.18U PW=1.18U
XI3 NET15 NET29 NET17 B TG1G NW=1.18U PW=1.18U
XI4 NET21 NET6 NET35 C TG1G NW=1.18U PW=1.18U
XI2 NET29 NET6 C NET35 TG1G NW=1.18U PW=1.18U
XI10 NET35 C IVG PW=0.64U NW=0.42U
XI7 NET13 A IVG PW=1.72U NW=1.22U
XI6 NET15 NET13 IVG PW=1.68U NW=1.18U
XI0 NET17 B IVG PW=0.96U NW=0.64U
XI1 Z NET6 IVG PW=2.4U NW=1.6U
.ENDS XOR3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR2HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:45:38 2002                                       *
*******************************************************************************
.SUBCKT XOR2HDLX Z A B
XI4 NET17 NET6 A NET19 TG1G NW=0.42U PW=0.42U
XI2 NET15 NET6 NET19 A TG1G NW=0.42U PW=0.42U
XI8 Z NET6 IVG PW=0.64U NW=0.42U
XI7 NET15 B IVG PW=0.45U NW=0.3U
XI6 NET17 NET15 IVG PW=0.45U NW=0.3U
XI0 NET19 A IVG PW=0.45U NW=0.3U
.ENDS XOR2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR2HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:45:30 2002                                       *
*******************************************************************************
.SUBCKT XOR2HD4X Z A B
XI2 NET11 NET18 NET7 A TG1G NW=2.44U PW=2.5U
XI3 NET9 NET18 A NET7 TG1G NW=2.44U PW=2.5U
XI1 Z NET18 IVG PW=4.8U NW=3.2U
XI0 NET7 A IVG PW=1.14U NW=0.76U
XI6 NET9 NET11 IVG PW=3.44U NW=2.4U
XI7 NET11 B IVG PW=6.48U NW=4.32U
.ENDS XOR2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR2HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:45:28 2002                                       *
*******************************************************************************
.SUBCKT XOR2HD2X Z A B
XI3 NET15 NET6 A NET17 TG1G NW=1.18U PW=1.2U
XI2 NET13 NET6 NET17 A TG1G NW=1.18U PW=1.2U
XI1 Z NET6 IVG PW=2.4U NW=1.6U
XI6 NET15 NET13 IVG PW=1.68U NW=1.18U
XI0 NET17 A IVG PW=0.64U NW=0.42U
XI7 NET13 B IVG PW=3.44U NW=2.32U
.ENDS XOR2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XOR2HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:45:26 2002                                       *
*******************************************************************************
.SUBCKT XOR2HD1X Z A B
XI4 NET19 NET6 A NET13 TG1G NW=0.6U PW=0.6U
XI2 NET17 NET6 NET13 A TG1G NW=0.6U PW=0.6U
XI8 Z NET6 IVG PW=1.2U NW=0.8U
XI7 NET17 B IVG PW=1.64U NW=1.12U
XI6 NET19 NET17 IVG PW=0.9U NW=0.6U
XI0 NET13 A IVG PW=0.45U NW=0.3U
.ENDS XOR2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR3HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:45:24 2002                                       *
*******************************************************************************
.SUBCKT XNOR3HD4X Z A B C
XI8 NET13 NET21 NET17 B TG1G NW=2U PW=2U
XI9 NET15 NET21 B NET17 TG1G NW=2U PW=2U
XI5 NET13 NET29 B NET17 TG1G NW=2U PW=2U
XI3 NET15 NET29 NET17 B TG1G NW=2U PW=2U
XI4 NET21 NET6 C NET35 TG1G NW=2U PW=2U
XI2 NET29 NET6 NET35 C TG1G NW=2U PW=2U
XI10 NET35 C IVG PW=0.9U NW=0.6U
XI7 NET13 A IVG PW=3.44U NW=2.4U
XI6 NET15 NET13 IVG PW=3.44U NW=2.4U
XI0 NET17 B IVG PW=1.68U NW=1.18U
XI1 Z NET6 IVG PW=4.8U NW=3.2U
.ENDS XNOR3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR3HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:45:22 2002                                       *
*******************************************************************************
.SUBCKT XNOR3HD2X Z A B C
XI8 NET13 NET21 NET17 B TG1G NW=1.18U PW=1.18U
XI9 NET15 NET21 B NET17 TG1G NW=1.18U PW=1.18U
XI5 NET13 NET29 B NET17 TG1G NW=1.18U PW=1.18U
XI3 NET15 NET29 NET17 B TG1G NW=1.18U PW=1.18U
XI4 NET21 NET6 C NET35 TG1G NW=1.18U PW=1.18U
XI2 NET29 NET6 NET35 C TG1G NW=1.18U PW=1.18U
XI10 NET35 C IVG PW=0.64U NW=0.42U
XI7 NET13 A IVG PW=1.72U NW=1.22U
XI6 NET15 NET13 IVG PW=1.68U NW=1.18U
XI0 NET17 B IVG PW=0.96U NW=0.64U
XI1 Z NET6 IVG PW=2.4U NW=1.6U
.ENDS XNOR3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR2HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:45:20 2002                                       *
*******************************************************************************
.SUBCKT XNOR2HDLX Z A B
XI0 NET5 A IVG PW=0.45U NW=0.3U
XI6 NET7 NET9 IVG PW=0.45U NW=0.3U
XI7 NET9 B IVG PW=0.45U NW=0.3U
XI8 Z NET18 IVG PW=0.64U NW=0.42U
XI2 NET9 NET18 A NET5 TG1G NW=0.42U PW=0.42U
XI4 NET7 NET18 NET5 A TG1G NW=0.42U PW=0.42U
.ENDS XNOR2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR2HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:45:18 2002                                       *
*******************************************************************************
.SUBCKT XNOR2HD4X Z A B
XI4 NET15 NET6 NET17 A TG1G NW=2.44U PW=2.5U
XI2 NET13 NET6 A NET17 TG1G NW=2.44U PW=2.5U
XI7 NET13 B IVG PW=6.48U NW=4.32U
XI6 NET15 NET13 IVG PW=3.44U NW=2.4U
XI0 NET17 A IVG PW=1.14U NW=0.76U
XI1 Z NET6 IVG PW=4.8U NW=3.2U
.ENDS XNOR2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR2HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:45:17 2002                                       *
*******************************************************************************
.SUBCKT XNOR2HD2X Z A B
XI1 Z NET18 IVG PW=2.4U NW=1.6U
XI0 NET7 A IVG PW=0.64U NW=0.42U
XI6 NET9 NET11 IVG PW=1.68U NW=1.18U
XI7 NET11 B IVG PW=3.44U NW=2.32U
XI2 NET11 NET18 A NET7 TG1G NW=1.18U PW=1.2U
XI4 NET9 NET18 NET7 A TG1G NW=1.18U PW=1.2U
.ENDS XNOR2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XNOR2HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:45:15 2002                                       *
*******************************************************************************
.SUBCKT XNOR2HD1X Z A B
XI4 NET15 NET19 NET17 A TG1G NW=0.6U PW=0.6U
XI2 NET13 NET19 A NET17 TG1G NW=0.6U PW=0.6U
XI8 Z NET19 IVG PW=1.2U NW=0.8U
XI7 NET13 B IVG PW=1.64U NW=1.12U
XI6 NET15 NET13 IVG PW=0.9U NW=0.6U
XI0 NET17 A IVG PW=0.45U NW=0.3U
.ENDS XNOR2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TIELHD                                                               *
* LAST TIME SAVED: AUG 30 10:44:06 2002                                       *
*******************************************************************************
.SUBCKT TIELHD Z
MP1 VDD NET5 NET5 VDD P18 W=0.3U L=0.18U
MN1 Z NET5 GND GND N18 W=0.56U L=0.18U
.ENDS TIELHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TIEHHD                                                               *
* LAST TIME SAVED: AUG 30 10:43:47 2002                                       *
*******************************************************************************
.SUBCKT TIEHHD Z
MN1 NET14 NET14 GND GND N18 W=0.42U L=0.18U
MP1 VDD NET14 Z VDD P18 W=1.2U L=0.18U
.ENDS TIEHHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NR2G                                                                 *
* LAST TIME SAVED: SEP 28 13:10:43 2001                                       *
*******************************************************************************
.SUBCKT NR2G Z A B PL=0.18U PW=0.24U NL=0.18U NW=0.24U
MN0 Z B GND GND N18 W=NW L=NL
MN2 Z A GND GND N18 W=NW L=NL
MP0 NET21 B Z VDD P18 W=PW L=PL
MP2 VDD A NET21 VDD P18 W=PW L=PL
.ENDS NR2G


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATNHDLX                                                           *
* LAST TIME SAVED: AUG 30 10:40:09 2002                                       *
*******************************************************************************
.SUBCKT RSLATNHDLX Q QN RN SN
XI18 NET9 NET49 NET43 NR2G PW=0.84U NW=0.42U
XI17 NET49 NET45 NET9 NR2G PW=0.84U NW=0.42U
XI19 Q NET9 IVG PW=0.64U NW=0.42U
XI20 NET45 RN IVG PW=0.64U NW=0.42U
XI22 NET43 SN IVG PW=0.64U NW=0.42U
XI5 QN NET49 IVG PW=0.64U NW=0.42U
.ENDS RSLATNHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATNHD4X                                                           *
* LAST TIME SAVED: AUG 30 10:40:07 2002                                       *
*******************************************************************************
.SUBCKT RSLATNHD4X Q QN RN SN
XI18 NET9 NET49 NET43 NR2G PW=3.36U NW=1.68U
XI17 NET49 NET45 NET9 NR2G PW=3.36U NW=1.68U
XI19 Q NET9 IVG PW=4.8U NW=3.2U
XI20 NET45 RN IVG PW=1.5U NW=1U
XI22 NET43 SN IVG PW=1.5U NW=1U
XI5 QN NET49 IVG PW=4.8U NW=3.2U
.ENDS RSLATNHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATNHD2X                                                           *
* LAST TIME SAVED: AUG 30 10:40:05 2002                                       *
*******************************************************************************
.SUBCKT RSLATNHD2X Q QN RN SN
XI18 NET9 NET49 NET43 NR2G PW=1.68U NW=0.84U
XI17 NET49 NET45 NET9 NR2G PW=1.68U NW=0.84U
XI19 Q NET9 IVG PW=2.4U NW=1.6U
XI20 NET45 RN IVG PW=0.75U NW=0.5U
XI22 NET43 SN IVG PW=0.75U NW=0.5U
XI5 QN NET49 IVG PW=2.4U NW=1.6U
.ENDS RSLATNHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATNHD1X                                                           *
* LAST TIME SAVED: AUG 30 10:40:03 2002                                       *
*******************************************************************************
.SUBCKT RSLATNHD1X Q QN RN SN
XI18 NET9 NET49 NET43 NR2G PW=1.2U NW=0.6U
XI17 NET49 NET45 NET9 NR2G PW=1.2U NW=0.6U
XI19 Q NET9 IVG PW=1.2U NW=0.8U
XI20 NET45 RN IVG PW=0.64U NW=0.42U
XI22 NET43 SN IVG PW=0.64U NW=0.42U
XI5 QN NET49 IVG PW=1.2U NW=0.8U
.ENDS RSLATNHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: ND2G                                                                 *
* LAST TIME SAVED: SEP 28 11:59:32 2001                                       *
*******************************************************************************
.SUBCKT ND2G Z A B PL=0.18U PW=0.24U NL=0.18U NW=0.24U
MN2 NET15 A GND GND N18 W=NW L=NL
MN0 Z B NET15 GND N18 W=NW L=NL
MP2 VDD A Z VDD P18 W=PW L=PL
MP0 VDD B Z VDD P18 W=PW L=PL
.ENDS ND2G


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATHDLX                                                            *
* LAST TIME SAVED: AUG 30 10:40:17 2002                                       *
*******************************************************************************
.SUBCKT RSLATHDLX Q QN R S
XI19 QN NET9 IVG PW=0.64U NW=0.42U
XI20 NET45 R IVG PW=0.64U NW=0.42U
XI22 NET43 S IVG PW=0.64U NW=0.42U
XI5 Q NET49 IVG PW=0.64U NW=0.42U
XI18 NET9 NET49 NET43 ND2G PW=0.51U NW=0.42U
XI17 NET49 NET45 NET9 ND2G PW=0.51U NW=0.42U
.ENDS RSLATHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATHD4X                                                            *
* LAST TIME SAVED: AUG 30 10:40:15 2002                                       *
*******************************************************************************
.SUBCKT RSLATHD4X Q QN R S
XI18 NET9 NET49 NET43 ND2G PW=2.84U NW=2.36U
XI17 NET49 NET45 NET9 ND2G PW=2.84U NW=2.36U
XI19 QN NET9 IVG PW=4.8U NW=3.2U
XI20 NET45 R IVG PW=1.56U NW=1.04U
XI22 NET43 S IVG PW=1.56U NW=1.04U
XI5 Q NET49 IVG PW=4.8U NW=3.2U
.ENDS RSLATHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATHD2X                                                            *
* LAST TIME SAVED: AUG 30 10:40:14 2002                                       *
*******************************************************************************
.SUBCKT RSLATHD2X Q QN R S
XI19 QN NET9 IVG PW=2.4U NW=1.6U
XI20 NET45 R IVG PW=0.78U NW=0.52U
XI22 NET43 S IVG PW=0.78U NW=0.52U
XI5 Q NET49 IVG PW=2.4U NW=1.6U
XI18 NET9 NET49 NET43 ND2G PW=1.42U NW=1.18U
XI17 NET49 NET45 NET9 ND2G PW=1.42U NW=1.18U
.ENDS RSLATHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: RSLATHD1X                                                            *
* LAST TIME SAVED: AUG 30 10:40:11 2002                                       *
*******************************************************************************
.SUBCKT RSLATHD1X Q QN R S
XI19 QN NET9 IVG PW=1.2U NW=0.8U
XI20 NET45 R IVG PW=0.64U NW=0.42U
XI22 NET43 S IVG PW=0.64U NW=0.42U
XI5 Q NET49 IVG PW=1.2U NW=0.8U
XI18 NET9 NET49 NET43 ND2G PW=0.96U NW=0.8U
XI17 NET49 NET45 NET9 ND2G PW=0.96U NW=0.8U
.ENDS RSLATHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PULLUHD                                                              *
* LAST TIME SAVED: AUG 30 10:40:01 2002                                       *
*******************************************************************************
.SUBCKT PULLUHD Z E
MN0 NET8 E GND GND N18 W=0.42U L=0.18U
MN1 VDD NET8 Z VDD P18 W=1.2U L=0.18U
MP0 VDD E NET8 VDD P18 W=0.64U L=0.18U
.ENDS PULLUHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PULLDHD                                                              *
* LAST TIME SAVED: AUG 30 10:40:00 2002                                       *
*******************************************************************************
.SUBCKT PULLDHD Z EN
MN1 Z NET8 GND GND N18 W=0.8U L=0.18U
MN0 NET8 EN GND GND N18 W=0.42U L=0.18U
MP0 VDD EN NET8 VDD P18 W=0.64U L=0.18U
.ENDS PULLDHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR4HDLX                                                              *
* LAST TIME SAVED: AUG 30 10:39:58 2002                                       *
*******************************************************************************
.SUBCKT OR4HDLX Z A B C D
XI4 Z NET25 IVG PW=0.64U NW=0.42U
MN4 NET25 A GND GND N18 W=0.42U L=0.18U
MN3 NET25 B GND GND N18 W=0.42U L=0.18U
MN2 NET25 D GND GND N18 W=0.42U L=0.18U
MN0 NET25 C GND GND N18 W=0.42U L=0.18U
MP4 NET38 D NET25 VDD P18 W=1.16U L=0.18U
MP3 NET27 C NET38 VDD P18 W=1.16U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.16U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.16U L=0.18U
.ENDS OR4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR4HD4X                                                              *
* LAST TIME SAVED: AUG 30 10:39:56 2002                                       *
*******************************************************************************
.SUBCKT OR4HD4X Z A B C D
XI4 Z NET25 IVG PW=4.8U NW=3.2U
MN4 NET25 A GND GND N18 W=0.6U L=0.18U
MN3 NET25 B GND GND N18 W=0.6U L=0.18U
MN2 NET25 D GND GND N18 W=0.6U L=0.18U
MN0 NET25 C GND GND N18 W=0.6U L=0.18U
MP4 NET38 D NET25 VDD P18 W=1.68U L=0.18U
MP3 NET27 C NET38 VDD P18 W=1.68U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
.ENDS OR4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR4HD2X                                                              *
* LAST TIME SAVED: AUG 30 10:39:55 2002                                       *
*******************************************************************************
.SUBCKT OR4HD2X Z A B C D
XI4 Z NET25 IVG PW=2.4U NW=1.6U
MN4 NET25 A GND GND N18 W=0.54U L=0.18U
MN3 NET25 B GND GND N18 W=0.54U L=0.18U
MN2 NET25 D GND GND N18 W=0.54U L=0.18U
MN0 NET25 C GND GND N18 W=0.54U L=0.18U
MP4 NET38 D NET25 VDD P18 W=1.48U L=0.18U
MP3 NET27 C NET38 VDD P18 W=1.48U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.48U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.48U L=0.18U
.ENDS OR4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR4HD1X                                                              *
* LAST TIME SAVED: AUG 30 10:39:53 2002                                       *
*******************************************************************************
.SUBCKT OR4HD1X Z A B C D
XI4 Z NET25 IVG PW=1.2U NW=0.8U
MN4 NET25 A GND GND N18 W=0.42U L=0.18U
MN3 NET25 B GND GND N18 W=0.42U L=0.18U
MN2 NET25 D GND GND N18 W=0.42U L=0.18U
MN0 NET25 C GND GND N18 W=0.42U L=0.18U
MP4 NET38 D NET25 VDD P18 W=1.16U L=0.18U
MP3 NET27 C NET38 VDD P18 W=1.16U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.16U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.16U L=0.18U
.ENDS OR4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR3HDLX                                                              *
* LAST TIME SAVED: AUG 30 10:39:51 2002                                       *
*******************************************************************************
.SUBCKT OR3HDLX Z A B C
XI4 Z NET22 IVG PW=0.64U NW=0.42U
MN3 NET22 A GND GND N18 W=0.42U L=0.18U
MN2 NET22 C GND GND N18 W=0.42U L=0.18U
MN0 NET22 B GND GND N18 W=0.42U L=0.18U
MP3 NET27 C NET22 VDD P18 W=1.0U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.0U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.0U L=0.18U
.ENDS OR3HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR3HD4X                                                              *
* LAST TIME SAVED: AUG 30 10:39:49 2002                                       *
*******************************************************************************
.SUBCKT OR3HD4X Z A B C
XI4 Z NET22 IVG PW=4.8U NW=3.2U
MN3 NET22 A GND GND N18 W=0.7U L=0.18U
MN2 NET22 C GND GND N18 W=0.7U L=0.18U
MN0 NET22 B GND GND N18 W=0.7U L=0.18U
MP3 NET27 C NET22 VDD P18 W=1.68U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
.ENDS OR3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR3HD2X                                                              *
* LAST TIME SAVED: AUG 30 10:39:47 2002                                       *
*******************************************************************************
.SUBCKT OR3HD2X Z A B C
XI4 Z NET22 IVG PW=2.4U NW=1.6U
MN3 NET22 A GND GND N18 W=0.54U L=0.18U
MN2 NET22 C GND GND N18 W=0.54U L=0.18U
MN0 NET22 B GND GND N18 W=0.54U L=0.18U
MP3 NET27 C NET22 VDD P18 W=1.3U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.3U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.3U L=0.18U
.ENDS OR3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR3HD1X                                                              *
* LAST TIME SAVED: AUG 30 10:39:46 2002                                       *
*******************************************************************************
.SUBCKT OR3HD1X Z A B C
XI4 Z NET22 IVG PW=1.2U NW=0.8U
MN3 NET22 A GND GND N18 W=0.42U L=0.18U
MN2 NET22 C GND GND N18 W=0.42U L=0.18U
MN0 NET22 B GND GND N18 W=0.42U L=0.18U
MP3 NET27 C NET22 VDD P18 W=1.0U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.0U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.0U L=0.18U
.ENDS OR3HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2ODHD                                                              *
* LAST TIME SAVED: AUG 30 10:39:33 2002                                       *
*******************************************************************************
.SUBCKT OR2ODHD Z A B
MP4 NET21 B NET9 VDD P18 W=1.6U L=0.18U
MP1 VDD A NET21 VDD P18 W=1.6U L=0.18U
MN2 Z NET9 GND GND N18 W=1.18U L=0.18U M=2
MN3 NET9 A GND GND N18 W=0.8U L=0.18U
MN4 NET9 B GND GND N18 W=0.8U L=0.18U
.ENDS OR2ODHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HDLX                                                              *
* LAST TIME SAVED: AUG 30 10:39:44 2002                                       *
*******************************************************************************
.SUBCKT OR2HDLX Z A B
XI4 Z NET21 IVG PW=0.64U NW=0.42U
MN2 NET21 B GND GND N18 W=0.42U L=0.18U
MN0 NET21 A GND GND N18 W=0.42U L=0.18U
MP1 VDD A NET12 VDD P18 W=0.84U L=0.18U
MP2 NET12 B NET21 VDD P18 W=0.84U L=0.18U
.ENDS OR2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HD4XSPG                                                           *
* LAST TIME SAVED: AUG 30 10:39:41 2002                                       *
*******************************************************************************
.SUBCKT OR2HD4XSPG Z A B
XI4 Z NET21 IVG PW=4.8U NW=3.2U
MN2 NET21 B GND GND N18 W=0.84U L=0.18U
MN0 NET21 A GND GND N18 W=0.84U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET21 VDD P18 W=1.68U L=0.18U
.ENDS OR2HD4XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HD4X                                                              *
* LAST TIME SAVED: AUG 30 10:39:40 2002                                       *
*******************************************************************************
.SUBCKT OR2HD4X Z A B
XI4 Z NET21 IVG PW=4.8U NW=3.2U
MN2 NET21 B GND GND N18 W=0.84U L=0.18U
MN0 NET21 A GND GND N18 W=0.84U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET21 VDD P18 W=1.68U L=0.18U
.ENDS OR2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HD2XSPG                                                           *
* LAST TIME SAVED: AUG 30 10:39:38 2002                                       *
*******************************************************************************
.SUBCKT OR2HD2XSPG Z A B
XI4 Z NET21 IVG PW=2.4U NW=1.6U
MN2 NET21 B GND GND N18 W=0.54U L=0.18U
MN0 NET21 A GND GND N18 W=0.54U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.08U L=0.18U
MP2 NET12 B NET21 VDD P18 W=1.08U L=0.18U
.ENDS OR2HD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HD2X                                                              *
* LAST TIME SAVED: AUG 30 10:39:36 2002                                       *
*******************************************************************************
.SUBCKT OR2HD2X Z A B
XI4 Z NET21 IVG PW=2.4U NW=1.6U
MN2 NET21 B GND GND N18 W=0.54U L=0.18U
MN0 NET21 A GND GND N18 W=0.54U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.08U L=0.18U
MP2 NET12 B NET21 VDD P18 W=1.08U L=0.18U
.ENDS OR2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OR2HD1X                                                              *
* LAST TIME SAVED: AUG 30 10:39:35 2002                                       *
*******************************************************************************
.SUBCKT OR2HD1X Z A B
XI4 Z NET21 IVG PW=1.2U NW=0.8U
MN2 NET21 B GND GND N18 W=0.42U L=0.18U
MN0 NET21 A GND GND N18 W=0.42U L=0.18U
MP1 VDD A NET12 VDD P18 W=0.84U L=0.18U
MP2 NET12 B NET21 VDD P18 W=0.84U L=0.18U
.ENDS OR2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI33HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:39:31 2002                                       *
*******************************************************************************
.SUBCKT OAI33HDLX Z A B C D E F
MP7 NET55 E NET40 VDD P18 W=1.0U L=0.18U
MP8 NET37 B NET12 VDD P18 W=1.0U L=0.18U
MP6 VDD F NET55 VDD P18 W=1.0U L=0.18U
MP9 NET40 D Z VDD P18 W=1.0U L=0.18U
MP2 VDD A NET37 VDD P18 W=1.0U L=0.18U
MP10 NET12 C Z VDD P18 W=1.0U L=0.18U
MN11 Z E NET64 GND N18 W=0.52U L=0.18U
MN12 Z D NET64 GND N18 W=0.52U L=0.18U
MN9 NET64 A GND GND N18 W=0.52U L=0.18U
MN8 NET64 B GND GND N18 W=0.52U L=0.18U
MN10 Z F NET64 GND N18 W=0.52U L=0.18U
MN0 NET64 C GND GND N18 W=0.52U L=0.18U
.ENDS OAI33HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI33HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:39:30 2002                                       *
*******************************************************************************
.SUBCKT OAI33HD4X Z A B C D E F
XI4 NET39 NET72 IVG PW=1.6U NW=1.06U
XI5 Z NET39 IVG PW=4.8U NW=3.2U
MP7 NET55 E NET40 VDD P18 W=1.0U L=0.18U
MP8 NET37 B NET12 VDD P18 W=1.0U L=0.18U
MP6 VDD F NET55 VDD P18 W=1.0U L=0.18U
MP9 NET40 D NET72 VDD P18 W=1.0U L=0.18U
MP2 VDD A NET37 VDD P18 W=1.0U L=0.18U
MP10 NET12 C NET72 VDD P18 W=1.0U L=0.18U
MN11 NET72 E NET64 GND N18 W=0.52U L=0.18U
MN12 NET72 D NET64 GND N18 W=0.52U L=0.18U
MN9 NET64 A GND GND N18 W=0.52U L=0.18U
MN8 NET64 B GND GND N18 W=0.52U L=0.18U
MN10 NET72 F NET64 GND N18 W=0.52U L=0.18U
MN0 NET64 C GND GND N18 W=0.52U L=0.18U
.ENDS OAI33HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI33HD2X                                                            *
* LAST TIME SAVED: JUL 14 11:31:04 2004                                       *
*******************************************************************************
.SUBCKT OAI33HD2X Z A B C D E F
XI4 NET39 NET72 IVG PW=0.8U NW=0.53U
XI5 Z NET39 IVG PW=2.4U NW=1.6U
MP7 NET55 E NET40 VDD P18 W=0.81U L=0.18U
MP8 NET37 B NET12 VDD P18 W=0.81U L=0.18U
MP6 VDD F NET55 VDD P18 W=0.81U L=0.18U
MP9 NET40 D NET72 VDD P18 W=0.81U L=0.18U
MP2 VDD A NET37 VDD P18 W=0.81U L=0.18U
MP10 NET12 C NET72 VDD P18 W=0.81U L=0.18U
MN11 NET72 E NET64 GND N18 W=0.42U L=0.18U
MN12 NET72 D NET64 GND N18 W=0.42U L=0.18U
MN9 NET64 A GND GND N18 W=0.42U L=0.18U
MN8 NET64 B GND GND N18 W=0.42U L=0.18U
MN10 NET72 F NET64 GND N18 W=0.42U L=0.18U
MN0 NET64 C GND GND N18 W=0.42U L=0.18U
.ENDS OAI33HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI33HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:39:26 2002                                       *
*******************************************************************************
.SUBCKT OAI33HD1X Z A B C D E F
MP7 NET55 E NET40 VDD P18 W=1.68U L=0.18U
MP8 NET37 B NET12 VDD P18 W=1.68U L=0.18U
MP6 VDD F NET55 VDD P18 W=1.68U L=0.18U
MP9 NET40 D Z VDD P18 W=1.68U L=0.18U
MP2 VDD A NET37 VDD P18 W=1.68U L=0.18U
MP10 NET12 C Z VDD P18 W=1.68U L=0.18U
MN11 Z E NET64 GND N18 W=0.88U L=0.18U
MN12 Z D NET64 GND N18 W=0.88U L=0.18U
MN9 NET64 A GND GND N18 W=0.88U L=0.18U
MN8 NET64 B GND GND N18 W=0.88U L=0.18U
MN10 Z F NET64 GND N18 W=0.88U L=0.18U
MN0 NET64 C GND GND N18 W=0.88U L=0.18U
.ENDS OAI33HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI32HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:39:25 2002                                       *
*******************************************************************************
.SUBCKT OAI32HDLX Z A B C D E
MP8 NET12 C Z VDD P18 W=1.0U L=0.18U
MP5 NET28 B NET12 VDD P18 W=1.0U L=0.18U
MP7 NET45 E Z VDD P18 W=0.84U L=0.18U
MP2 VDD A NET28 VDD P18 W=1.0U L=0.18U
MP6 VDD D NET45 VDD P18 W=0.84U L=0.18U
MN7 NET37 B GND GND N18 W=0.52U L=0.18U
MN8 NET37 C GND GND N18 W=0.52U L=0.18U
MN9 Z E NET37 GND N18 W=0.52U L=0.18U
MN10 Z D NET37 GND N18 W=0.52U L=0.18U
MN5 NET37 A GND GND N18 W=0.52U L=0.18U
.ENDS OAI32HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI32HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:39:23 2002                                       *
*******************************************************************************
.SUBCKT OAI32HD4X Z A B C D E
XI4 NET34 NET64 IVG PW=1.6U NW=1.06U
XI5 Z NET34 IVG PW=4.8U NW=3.2U
MP8 NET12 C NET64 VDD P18 W=1.0U L=0.18U
MP5 NET28 B NET12 VDD P18 W=1.0U L=0.18U
MP7 NET45 E NET64 VDD P18 W=0.84U L=0.18U
MP2 VDD A NET28 VDD P18 W=1.0U L=0.18U
MP6 VDD D NET45 VDD P18 W=0.84U L=0.18U
MN7 NET37 B GND GND N18 W=0.52U L=0.18U
MN8 NET37 C GND GND N18 W=0.52U L=0.18U
MN9 NET64 E NET37 GND N18 W=0.52U L=0.18U
MN10 NET64 D NET37 GND N18 W=0.52U L=0.18U
MN5 NET37 A GND GND N18 W=0.52U L=0.18U
.ENDS OAI32HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI32HD2X                                                            *
* LAST TIME SAVED: JUL 14 11:29:13 2004                                       *
*******************************************************************************
.SUBCKT OAI32HD2X Z A B C D E
XI4 NET34 NET64 IVG PW=0.8U NW=0.53U
XI5 Z NET34 IVG PW=2.4U NW=1.6U
MP8 NET12 C NET64 VDD P18 W=0.81U L=0.18U
MP5 NET28 B NET12 VDD P18 W=0.81U L=0.18U
MP7 NET45 E NET64 VDD P18 W=0.68U L=0.18U
MP2 VDD A NET28 VDD P18 W=0.81U L=0.18U
MP6 VDD D NET45 VDD P18 W=0.68U L=0.18U
MN7 NET37 B GND GND N18 W=0.42U L=0.18U
MN8 NET37 C GND GND N18 W=0.42U L=0.18U
MN9 NET64 E NET37 GND N18 W=0.42U L=0.18U
MN10 NET64 D NET37 GND N18 W=0.42U L=0.18U
MN5 NET37 A GND GND N18 W=0.42U L=0.18U
.ENDS OAI32HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI32HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:39:20 2002                                       *
*******************************************************************************
.SUBCKT OAI32HD1X Z A B C D E
MP8 NET12 C Z VDD P18 W=1.68U L=0.18U
MP5 NET28 B NET12 VDD P18 W=1.68U L=0.18U
MP7 NET45 E Z VDD P18 W=1.6U L=0.18U
MP2 VDD A NET28 VDD P18 W=1.68U L=0.18U
MP6 VDD D NET45 VDD P18 W=1.6U L=0.18U
MN7 NET37 B GND GND N18 W=0.88U L=0.18U
MN8 NET37 C GND GND N18 W=0.88U L=0.18U
MN9 Z E NET37 GND N18 W=1.0U L=0.18U
MN10 Z D NET37 GND N18 W=1.0U L=0.18U
MN5 NET37 A GND GND N18 W=0.88U L=0.18U
.ENDS OAI32HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI31HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:39:19 2002                                       *
*******************************************************************************
.SUBCKT OAI31HDLX Z A B C D
MP5 NET12 C Z VDD P18 W=1.0U L=0.18U
MP2 VDD A NET35 VDD P18 W=1.0U L=0.18U
MP6 VDD D Z VDD P18 W=0.64U L=0.18U
MP4 NET35 B NET12 VDD P18 W=1.0U L=0.18U
MN7 NET37 A GND GND N18 W=0.52U L=0.18U
MN8 Z D NET37 GND N18 W=0.52U L=0.18U
MN6 NET37 B GND GND N18 W=0.52U L=0.18U
MN5 NET37 C GND GND N18 W=0.52U L=0.18U
.ENDS OAI31HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI31HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:39:17 2002                                       *
*******************************************************************************
.SUBCKT OAI31HD4X Z A B C D
XI4 NET27 NET38 IVG PW=1.6U NW=1.06U
XI5 Z NET27 IVG PW=4.8U NW=3.2U
MP5 NET12 C NET38 VDD P18 W=1.0U L=0.18U
MP2 VDD A NET35 VDD P18 W=1.0U L=0.18U
MP6 VDD D NET38 VDD P18 W=0.64U L=0.18U
MP4 NET35 B NET12 VDD P18 W=1.0U L=0.18U
MN7 NET37 A GND GND N18 W=0.52U L=0.18U
MN8 NET38 D NET37 GND N18 W=0.52U L=0.18U
MN6 NET37 B GND GND N18 W=0.52U L=0.18U
MN5 NET37 C GND GND N18 W=0.52U L=0.18U
.ENDS OAI31HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI31HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:39:15 2002                                       *
*******************************************************************************
.SUBCKT OAI31HD2X Z A B C D
MP5 NET12 C Z VDD P18 W=3.36U L=0.18U
MP2 VDD A NET35 VDD P18 W=3.36U L=0.18U
MP6 VDD D Z VDD P18 W=2.4U L=0.18U
MP4 NET35 B NET12 VDD P18 W=3.36U L=0.18U
MN7 NET37 A GND GND N18 W=1.76U L=0.18U
MN8 Z D NET37 GND N18 W=2.0U L=0.18U
MN6 NET37 B GND GND N18 W=1.76U L=0.18U
MN5 NET37 C GND GND N18 W=1.76U L=0.18U
.ENDS OAI31HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI31HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:39:13 2002                                       *
*******************************************************************************
.SUBCKT OAI31HD1X Z A B C D
MP5 NET12 C Z VDD P18 W=1.68U L=0.18U
MP2 VDD A NET35 VDD P18 W=1.68U L=0.18U
MP6 VDD D Z VDD P18 W=1.2U L=0.18U
MP4 NET35 B NET12 VDD P18 W=1.68U L=0.18U
MN7 NET37 A GND GND N18 W=0.88U L=0.18U
MN8 Z D NET37 GND N18 W=1.0U L=0.18U
MN6 NET37 B GND GND N18 W=0.88U L=0.18U
MN5 NET37 C GND GND N18 W=0.88U L=0.18U
.ENDS OAI31HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:39:00 2002                                       *
*******************************************************************************
.SUBCKT OAI22HDLX Z A B C D
MP3 VDD A NET12 VDD P18 W=0.84U L=0.18U
MP4 NET29 D Z VDD P18 W=0.84U L=0.18U
MP5 NET12 B Z VDD P18 W=0.84U L=0.18U
MP6 VDD C NET29 VDD P18 W=0.84U L=0.18U
MN8 Z D NET8 GND N18 W=0.54U L=0.18U
MN6 NET8 A GND GND N18 W=0.54U L=0.18U
MN5 Z C NET8 GND N18 W=0.54U L=0.18U
MN7 NET8 B GND GND N18 W=0.54U L=0.18U
.ENDS OAI22HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:38:59 2002                                       *
*******************************************************************************
.SUBCKT OAI22HD4X Z A B C D
MP3 VDD A NET12 VDD P18 W=6.4U L=0.18U
MP4 NET29 D Z VDD P18 W=6.4U L=0.18U
MP5 NET12 B Z VDD P18 W=6.4U L=0.18U
MP6 VDD C NET29 VDD P18 W=6.4U L=0.18U
MN8 Z D NET8 GND N18 W=3.66U L=0.18U
MN6 NET8 A GND GND N18 W=3.66U L=0.18U
MN5 Z C NET8 GND N18 W=3.66U L=0.18U
MN7 NET8 B GND GND N18 W=3.66U L=0.18U
.ENDS OAI22HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:38:57 2002                                       *
*******************************************************************************
.SUBCKT OAI22HD2X Z A B C D
MP3 VDD A NET12 VDD P18 W=3.2U L=0.18U
MP4 NET29 D Z VDD P18 W=3.2U L=0.18U
MP5 NET12 B Z VDD P18 W=3.2U L=0.18U
MP6 VDD C NET29 VDD P18 W=3.2U L=0.18U
MN8 Z D NET8 GND N18 W=2.0U L=0.18U
MN6 NET8 A GND GND N18 W=2.0U L=0.18U
MN5 Z C NET8 GND N18 W=2.0U L=0.18U
MN7 NET8 B GND GND N18 W=2.0U L=0.18U
.ENDS OAI22HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:38:56 2002                                       *
*******************************************************************************
.SUBCKT OAI22HD1X Z A B C D
MP3 VDD A NET12 VDD P18 W=1.6U L=0.18U
MP4 NET29 D Z VDD P18 W=1.6U L=0.18U
MP5 NET12 B Z VDD P18 W=1.6U L=0.18U
MP6 VDD C NET29 VDD P18 W=1.6U L=0.18U
MN8 Z D NET8 GND N18 W=1.0U L=0.18U
MN6 NET8 A GND GND N18 W=1.0U L=0.18U
MN5 Z C NET8 GND N18 W=1.0U L=0.18U
MN7 NET8 B GND GND N18 W=1.0U L=0.18U
.ENDS OAI22HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22B2HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:39:12 2002                                       *
*******************************************************************************
.SUBCKT OAI22B2HDLX Z AN BN C D
MP7 NET12 D Z VDD P18 W=0.84U L=0.18U
MP9 VDD AN NET35 VDD P18 W=0.64U L=0.18U
MP5 VDD NET35 Z VDD P18 W=0.64U L=0.18U
MP8 VDD BN NET35 VDD P18 W=0.64U L=0.18U
MP4 VDD C NET12 VDD P18 W=0.84U L=0.18U
MN7 Z NET35 NET8 GND N18 W=0.54U L=0.18U
MN8 NET8 C GND GND N18 W=0.54U L=0.18U
MN9 NET8 D GND GND N18 W=0.54U L=0.18U
MN11 NET48 AN GND GND N18 W=0.54U L=0.18U
MN10 NET35 BN NET48 GND N18 W=0.54U L=0.18U
.ENDS OAI22B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22B2HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:39:11 2002                                       *
*******************************************************************************
.SUBCKT OAI22B2HD4X Z AN BN C D
MP7 NET12 D Z VDD P18 W=6.4U L=0.18U
MP9 VDD AN NET35 VDD P18 W=1.42U L=0.18U
MP5 VDD NET35 Z VDD P18 W=4.8U L=0.18U
MP8 VDD BN NET35 VDD P18 W=1.42U L=0.18U
MP4 VDD C NET12 VDD P18 W=6.4U L=0.18U
MN7 Z NET35 NET8 GND N18 W=3.66U L=0.18U
MN8 NET8 C GND GND N18 W=3.66U L=0.18U
MN9 NET8 D GND GND N18 W=3.66U L=0.18U
MN11 NET48 AN GND GND N18 W=1.18U L=0.18U
MN10 NET35 BN NET48 GND N18 W=1.18U L=0.18U
.ENDS OAI22B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22B2HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:39:08 2002                                       *
*******************************************************************************
.SUBCKT OAI22B2HD2X Z AN BN C D
MP7 NET12 D Z VDD P18 W=3.2U L=0.18U
MP9 VDD AN NET35 VDD P18 W=1.0U L=0.18U
MP5 VDD NET35 Z VDD P18 W=2.4U L=0.18U
MP8 VDD BN NET35 VDD P18 W=1.0U L=0.18U
MP4 VDD C NET12 VDD P18 W=3.2U L=0.18U
MN7 Z NET35 NET8 GND N18 W=2.0U L=0.18U
MN8 NET8 C GND GND N18 W=2.0U L=0.18U
MN9 NET8 D GND GND N18 W=2.0U L=0.18U
MN11 NET48 AN GND GND N18 W=0.84U L=0.18U
MN10 NET35 BN NET48 GND N18 W=0.84U L=0.18U
.ENDS OAI22B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI22B2HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:39:07 2002                                       *
*******************************************************************************
.SUBCKT OAI22B2HD1X Z AN BN C D
MP7 NET12 D Z VDD P18 W=1.6U L=0.18U
MP9 VDD AN NET35 VDD P18 W=0.64U L=0.18U
MP5 VDD NET35 Z VDD P18 W=1.2U L=0.18U
MP8 VDD BN NET35 VDD P18 W=0.64U L=0.18U
MP4 VDD C NET12 VDD P18 W=1.6U L=0.18U
MN7 Z NET35 NET8 GND N18 W=1.0U L=0.18U
MN8 NET8 C GND GND N18 W=1.0U L=0.18U
MN9 NET8 D GND GND N18 W=1.0U L=0.18U
MN11 NET48 AN GND GND N18 W=0.54U L=0.18U
MN10 NET35 BN NET48 GND N18 W=0.54U L=0.18U
.ENDS OAI22B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI222HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:38:54 2002                                       *
*******************************************************************************
.SUBCKT OAI222HDLX Z A B C D E F
MP11 Z B NET38 VDD P18 W=0.84U L=0.18U
MP10 Z D NET43 VDD P18 W=0.84U L=0.18U
MP9 Z F NET55 VDD P18 W=0.84U L=0.18U
MP8 NET55 E VDD VDD P18 W=0.84U L=0.18U
MP7 NET43 C VDD VDD P18 W=0.84U L=0.18U
MP0 NET38 A VDD VDD P18 W=0.84U L=0.18U
MN12 Z E NET25 GND N18 W=0.56U L=0.18U
MN9 NET25 C NET12 GND N18 W=0.56U L=0.18U
MN10 NET25 D NET12 GND N18 W=0.56U L=0.18U
MN4 NET12 B GND GND N18 W=0.56U L=0.18U
MN8 NET12 A GND GND N18 W=0.56U L=0.18U
MN11 Z F NET25 GND N18 W=0.56U L=0.18U
.ENDS OAI222HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI222HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:38:52 2002                                       *
*******************************************************************************
.SUBCKT OAI222HD4X Z A B C D E F
XI4 NET40 NET49 IVG PW=1.6U NW=1.06U
XI5 Z NET40 IVG PW=4.8U NW=3.2U
MP11 NET49 B NET38 VDD P18 W=0.84U L=0.18U
MP10 NET49 D NET43 VDD P18 W=0.84U L=0.18U
MP9 NET49 F NET55 VDD P18 W=0.84U L=0.18U
MP8 NET55 E VDD VDD P18 W=0.84U L=0.18U
MP7 NET43 C VDD VDD P18 W=0.84U L=0.18U
MP0 NET38 A VDD VDD P18 W=0.84U L=0.18U
MN12 NET49 E NET25 GND N18 W=0.56U L=0.18U
MN9 NET25 C NET12 GND N18 W=0.56U L=0.18U
MN10 NET25 D NET12 GND N18 W=0.56U L=0.18U
MN4 NET12 B GND GND N18 W=0.56U L=0.18U
MN8 NET12 A GND GND N18 W=0.56U L=0.18U
MN11 NET49 F NET25 GND N18 W=0.56U L=0.18U
.ENDS OAI222HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI222HD2X                                                           *
* LAST TIME SAVED: JUL 14 11:25:26 2004                                       *
*******************************************************************************
.SUBCKT OAI222HD2X Z A B C D E F
XI4 NET40 NET49 IVG PW=0.8U NW=0.53U
XI5 Z NET40 IVG PW=2.4U NW=1.6U
MP11 NET49 B NET38 VDD P18 W=0.64U L=0.18U
MP10 NET49 D NET43 VDD P18 W=0.64U L=0.18U
MP9 NET49 F NET55 VDD P18 W=0.64U L=0.18U
MP8 NET55 E VDD VDD P18 W=0.64U L=0.18U
MP7 NET43 C VDD VDD P18 W=0.64U L=0.18U
MP0 NET38 A VDD VDD P18 W=0.64U L=0.18U
MN12 NET49 E NET25 GND N18 W=0.42U L=0.18U
MN9 NET25 C NET12 GND N18 W=0.42U L=0.18U
MN10 NET25 D NET12 GND N18 W=0.42U L=0.18U
MN4 NET12 B GND GND N18 W=0.42U L=0.18U
MN8 NET12 A GND GND N18 W=0.42U L=0.18U
MN11 NET49 F NET25 GND N18 W=0.42U L=0.18U
.ENDS OAI222HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI222HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:38:49 2002                                       *
*******************************************************************************
.SUBCKT OAI222HD1X Z A B C D E F
MP11 Z B NET38 VDD P18 W=1.6U L=0.18U
MP10 Z D NET43 VDD P18 W=1.6U L=0.18U
MP9 Z F NET55 VDD P18 W=1.6U L=0.18U
MP8 NET55 E VDD VDD P18 W=1.6U L=0.18U
MP7 NET43 C VDD VDD P18 W=1.6U L=0.18U
MP0 NET38 A VDD VDD P18 W=1.6U L=0.18U
MN12 Z E NET25 GND N18 W=1.1U L=0.18U
MN9 NET25 C NET12 GND N18 W=1.1U L=0.18U
MN10 NET25 D NET12 GND N18 W=1.1U L=0.18U
MN4 NET12 B GND GND N18 W=1.1U L=0.18U
MN8 NET12 A GND GND N18 W=1.1U L=0.18U
MN11 Z F NET25 GND N18 W=1.1U L=0.18U
.ENDS OAI222HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI221HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:38:47 2002                                       *
*******************************************************************************
.SUBCKT OAI221HDLX Z A B C D E
MP9 NET12 B Z VDD P18 W=0.84U L=0.18U
MP6 VDD C NET43 VDD P18 W=0.84U L=0.18U
MP8 NET43 D Z VDD P18 W=0.84U L=0.18U
MP7 VDD E Z VDD P18 W=0.64U L=0.18U
MP0 VDD A NET12 VDD P18 W=0.84U L=0.18U
MN10 Z E NET25 GND N18 W=0.56U L=0.18U
MN9 NET25 D NET57 GND N18 W=0.56U L=0.18U
MN7 NET57 A GND GND N18 W=0.56U L=0.18U
MN8 NET25 C NET57 GND N18 W=0.56U L=0.18U
MN0 NET57 B GND GND N18 W=0.56U L=0.18U
.ENDS OAI221HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI221HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:38:45 2002                                       *
*******************************************************************************
.SUBCKT OAI221HD4X Z A B C D E
XI4 NET35 NET46 IVG PW=1.6U NW=1.06U
XI5 Z NET35 IVG PW=4.8U NW=3.2U
MP9 NET12 B NET46 VDD P18 W=0.84U L=0.18U
MP6 VDD C NET43 VDD P18 W=0.84U L=0.18U
MP8 NET43 D NET46 VDD P18 W=0.84U L=0.18U
MP7 VDD E NET46 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET12 VDD P18 W=0.84U L=0.18U
MN10 NET46 E NET25 GND N18 W=0.56U L=0.18U
MN9 NET25 D NET57 GND N18 W=0.56U L=0.18U
MN7 NET57 A GND GND N18 W=0.56U L=0.18U
MN8 NET25 C NET57 GND N18 W=0.56U L=0.18U
MN0 NET57 B GND GND N18 W=0.56U L=0.18U
.ENDS OAI221HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI221HD2X                                                           *
* LAST TIME SAVED: JUL 14 16:02:17 2004                                       *
*******************************************************************************
.SUBCKT OAI221HD2X Z A B C D E
XI4 NET35 NET46 IVG PW=0.8U NW=0.53U
XI5 Z NET35 IVG PW=2.4U NW=1.6U
MP9 NET12 B NET46 VDD P18 W=0.84U L=0.18U
MP6 VDD C NET43 VDD P18 W=0.84U L=0.18U
MP8 NET43 D NET46 VDD P18 W=0.84U L=0.18U
MP7 VDD E NET46 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET12 VDD P18 W=0.84U L=0.18U
MN10 NET46 E NET25 GND N18 W=0.56U L=0.18U
MN9 NET25 D NET57 GND N18 W=0.56U L=0.18U
MN7 NET57 A GND GND N18 W=0.56U L=0.18U
MN8 NET25 C NET57 GND N18 W=0.56U L=0.18U
MN0 NET57 B GND GND N18 W=0.56U L=0.18U
.ENDS OAI221HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI221HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:38:42 2002                                       *
*******************************************************************************
.SUBCKT OAI221HD1X Z A B C D E
MP9 NET12 B Z VDD P18 W=1.6U L=0.18U
MP6 VDD C NET43 VDD P18 W=1.6U L=0.18U
MP8 NET43 D Z VDD P18 W=1.6U L=0.18U
MP7 VDD E Z VDD P18 W=1.2U L=0.18U
MP0 VDD A NET12 VDD P18 W=1.6U L=0.18U
MN10 Z E NET25 GND N18 W=1.1U L=0.18U
MN9 NET25 D NET57 GND N18 W=1.1U L=0.18U
MN7 NET57 A GND GND N18 W=1.1U L=0.18U
MN8 NET25 C NET57 GND N18 W=1.1U L=0.18U
MN0 NET57 B GND GND N18 W=1.1U L=0.18U
.ENDS OAI221HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:38:40 2002                                       *
*******************************************************************************
.SUBCKT OAI21HDLX Z A B C
MP3 VDD A NET12 VDD P18 W=0.84U L=0.18U
MP4 VDD C Z VDD P18 W=0.64U L=0.18U
MP5 NET12 B Z VDD P18 W=0.84U L=0.18U
MN6 NET8 A GND GND N18 W=0.54U L=0.18U
MN5 Z C NET8 GND N18 W=0.54U L=0.18U
MN7 NET8 B GND GND N18 W=0.54U L=0.18U
.ENDS OAI21HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:38:38 2002                                       *
*******************************************************************************
.SUBCKT OAI21HD4X Z A B C
MP3 VDD A NET12 VDD P18 W=6.4U L=0.18U
MP4 VDD C Z VDD P18 W=4.8U L=0.18U
MP5 NET12 B Z VDD P18 W=6.4U L=0.18U
MN6 NET8 A GND GND N18 W=3.2U L=0.18U
MN5 Z C NET8 GND N18 W=3.66U L=0.18U
MN7 NET8 B GND GND N18 W=3.66U L=0.18U
.ENDS OAI21HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:38:35 2002                                       *
*******************************************************************************
.SUBCKT OAI21HD2X Z A B C
MP3 VDD A NET12 VDD P18 W=3.2U L=0.18U
MP4 VDD C Z VDD P18 W=2.4U L=0.18U
MP5 NET12 B Z VDD P18 W=3.2U L=0.18U
MN6 NET8 A GND GND N18 W=2.0U L=0.18U
MN5 Z C NET8 GND N18 W=2.0U L=0.18U
MN7 NET8 B GND GND N18 W=2.0U L=0.18U
.ENDS OAI21HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:38:34 2002                                       *
*******************************************************************************
.SUBCKT OAI21HD1X Z A B C
MP3 VDD A NET12 VDD P18 W=1.6U L=0.18U
MP4 VDD C Z VDD P18 W=1.2U L=0.18U
MP5 NET12 B Z VDD P18 W=1.6U L=0.18U
MN6 NET8 A GND GND N18 W=1.0U L=0.18U
MN5 Z C NET8 GND N18 W=1.0U L=0.18U
MN7 NET8 B GND GND N18 W=1.0U L=0.18U
.ENDS OAI21HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21B2HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:39:07 2002                                       *
*******************************************************************************
.SUBCKT OAI21B2HDLX Z AN BN C
MP7 VDD AN NET35 VDD P18 W=0.64U L=0.18U
MP8 VDD C Z VDD P18 W=0.64U L=0.18U
MP9 VDD NET35 Z VDD P18 W=0.64U L=0.18U
MP5 VDD BN NET35 VDD P18 W=0.64U L=0.18U
MN7 NET35 BN NET45 GND N18 W=0.54U L=0.18U
MN8 NET45 AN GND GND N18 W=0.54U L=0.18U
MN9 NET42 C GND GND N18 W=0.54U L=0.18U
MN10 Z NET35 NET42 GND N18 W=0.54U L=0.18U
.ENDS OAI21B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21B2HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:39:05 2002                                       *
*******************************************************************************
.SUBCKT OAI21B2HD4X Z AN BN C
MP7 VDD AN NET35 VDD P18 W=1.42U L=0.18U
MP8 VDD C Z VDD P18 W=4.8U L=0.18U
MP9 VDD NET35 Z VDD P18 W=4.8U L=0.18U
MP5 VDD BN NET35 VDD P18 W=1.42U L=0.18U
MN7 NET35 BN NET45 GND N18 W=1.18U L=0.18U
MN8 NET45 AN GND GND N18 W=1.18U L=0.18U
MN9 NET42 C GND GND N18 W=3.66U L=0.18U
MN10 Z NET35 NET42 GND N18 W=3.66U L=0.18U
.ENDS OAI21B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21B2HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:39:04 2002                                       *
*******************************************************************************
.SUBCKT OAI21B2HD2X Z AN BN C
MP7 VDD AN NET35 VDD P18 W=0.8U L=0.18U
MP8 VDD C Z VDD P18 W=2.4U L=0.18U
MP9 VDD NET35 Z VDD P18 W=2.4U L=0.18U
MP5 VDD BN NET35 VDD P18 W=0.8U L=0.18U
MN7 NET35 BN NET45 GND N18 W=0.64U L=0.18U
MN8 NET45 AN GND GND N18 W=0.64U L=0.18U
MN9 NET42 C GND GND N18 W=2.0U L=0.18U
MN10 Z NET35 NET42 GND N18 W=2.0U L=0.18U
.ENDS OAI21B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI21B2HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:39:02 2002                                       *
*******************************************************************************
.SUBCKT OAI21B2HD1X Z AN BN C
MP7 VDD AN NET35 VDD P18 W=0.64U L=0.18U
MP8 VDD C Z VDD P18 W=1.2U L=0.18U
MP9 VDD NET35 Z VDD P18 W=1.2U L=0.18U
MP5 VDD BN NET35 VDD P18 W=0.64U L=0.18U
MN7 NET35 BN NET45 GND N18 W=0.54U L=0.18U
MN8 NET45 AN GND GND N18 W=0.54U L=0.18U
MN9 NET42 C GND GND N18 W=1.0U L=0.18U
MN10 Z NET35 NET42 GND N18 W=1.0U L=0.18U
.ENDS OAI21B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI211HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:38:32 2002                                       *
*******************************************************************************
.SUBCKT OAI211HDLX Z A B C D
MP4 NET26 B Z VDD P18 W=0.84U L=0.18U
MP5 VDD D Z VDD P18 W=0.64U L=0.18U
MP3 VDD A NET26 VDD P18 W=0.84U L=0.18U
MP6 VDD C Z VDD P18 W=0.64U L=0.18U
MN6 NET12 A GND GND N18 W=0.58U L=0.18U
MN7 NET18 C NET12 GND N18 W=0.58U L=0.18U
MN8 Z D NET18 GND N18 W=0.58U L=0.18U
MN4 NET12 B GND GND N18 W=0.58U L=0.18U
.ENDS OAI211HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI211HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:38:30 2002                                       *
*******************************************************************************
.SUBCKT OAI211HD4X Z A B C D
XI4 NET54 NET39 IVG PW=1.6U NW=1.06U
XI5 Z NET54 IVG PW=4.8U NW=3.2U
MP4 NET26 B NET39 VDD P18 W=0.84U L=0.18U
MP5 VDD D NET39 VDD P18 W=0.64U L=0.18U
MP3 VDD A NET26 VDD P18 W=0.84U L=0.18U
MP6 VDD C NET39 VDD P18 W=0.64U L=0.18U
MN6 NET12 A GND GND N18 W=0.58U L=0.18U
MN7 NET18 C NET12 GND N18 W=0.58U L=0.18U
MN8 NET39 D NET18 GND N18 W=0.58U L=0.18U
MN4 NET12 B GND GND N18 W=0.58U L=0.18U
.ENDS OAI211HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI211HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:38:28 2002                                       *
*******************************************************************************
.SUBCKT OAI211HD2X Z A B C D
MP4 NET26 B Z VDD P18 W=3.2U L=0.18U
MP5 VDD D Z VDD P18 W=2.4U L=0.18U
MP3 VDD A NET26 VDD P18 W=3.2U L=0.18U
MP6 VDD C Z VDD P18 W=2.4U L=0.18U
MN6 NET12 A GND GND N18 W=2.2U L=0.18U
MN7 NET18 C NET12 GND N18 W=2.2U L=0.18U
MN8 Z D NET18 GND N18 W=2.2U L=0.18U
MN4 NET12 B GND GND N18 W=2.2U L=0.18U
.ENDS OAI211HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OAI211HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:38:28 2002                                       *
*******************************************************************************
.SUBCKT OAI211HD1X Z A B C D
MP4 NET26 B Z VDD P18 W=1.6U L=0.18U
MP5 VDD D Z VDD P18 W=1.2U L=0.18U
MP3 VDD A NET26 VDD P18 W=1.6U L=0.18U
MP6 VDD C Z VDD P18 W=1.2U L=0.18U
MN6 NET12 A GND GND N18 W=1.1U L=0.18U
MN7 NET18 C NET12 GND N18 W=1.1U L=0.18U
MN8 Z D NET18 GND N18 W=1.1U L=0.18U
MN4 NET12 B GND GND N18 W=1.1U L=0.18U
.ENDS OAI211HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:38:26 2002                                       *
*******************************************************************************
.SUBCKT NOR4HDLX Z A B C D
MN4 Z A GND GND N18 W=0.42U L=0.18U
MN3 Z B GND GND N18 W=0.42U L=0.18U
MN2 Z D GND GND N18 W=0.42U L=0.18U
MN0 Z C GND GND N18 W=0.42U L=0.18U
MP4 NET35 D Z VDD P18 W=1.16U L=0.18U
MP3 NET27 C NET35 VDD P18 W=1.16U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.16U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.16U L=0.18U
.ENDS NOR4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:38:24 2002                                       *
*******************************************************************************
.SUBCKT NOR4HD4X Z A B C D
MN4 Z A GND GND N18 W=2.4U L=0.18U
MN3 Z B GND GND N18 W=2.4U L=0.18U
MN2 Z D GND GND N18 W=2.4U L=0.18U
MN0 Z C GND GND N18 W=2.4U L=0.18U
MP4 NET35 D Z VDD P18 W=6.72U L=0.18U
MP3 NET27 C NET35 VDD P18 W=6.72U L=0.18U
MP1 VDD A NET12 VDD P18 W=6.72U L=0.18U
MP2 NET12 B NET27 VDD P18 W=6.72U L=0.18U
.ENDS NOR4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:38:23 2002                                       *
*******************************************************************************
.SUBCKT NOR4HD2X Z A B C D
MN4 Z A GND GND N18 W=1.2U L=0.18U
MN3 Z B GND GND N18 W=1.2U L=0.18U
MN2 Z D GND GND N18 W=1.2U L=0.18U
MN0 Z C GND GND N18 W=1.2U L=0.18U
MP4 NET35 D Z VDD P18 W=3.36U L=0.18U
MP3 NET27 C NET35 VDD P18 W=3.36U L=0.18U
MP1 VDD A NET12 VDD P18 W=3.36U L=0.18U
MP2 NET12 B NET27 VDD P18 W=3.36U L=0.18U
.ENDS NOR4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:38:21 2002                                       *
*******************************************************************************
.SUBCKT NOR4HD1X Z A B C D
MN4 Z A GND GND N18 W=0.6U L=0.18U
MN3 Z B GND GND N18 W=0.6U L=0.18U
MN2 Z D GND GND N18 W=0.6U L=0.18U
MN0 Z C GND GND N18 W=0.6U L=0.18U
MP4 NET35 D Z VDD P18 W=1.68U L=0.18U
MP3 NET27 C NET35 VDD P18 W=1.68U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
.ENDS NOR4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B2HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:38:12 2002                                       *
*******************************************************************************
.SUBCKT NOR4B2HDLX Z AN BN C D
MN4 Z NET17 GND GND N18 W=0.42U L=0.18U
MN3 Z NET47 GND GND N18 W=0.42U L=0.18U
MN2 Z D GND GND N18 W=0.42U L=0.18U
MN0 Z C GND GND N18 W=0.42U L=0.18U
MP4 NET37 D Z VDD P18 W=1.16U L=0.18U
MP3 NET27 C NET37 VDD P18 W=1.16U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.16U L=0.18U
MP2 NET12 NET47 NET27 VDD P18 W=1.16U L=0.18U
XI4 NET47 BN IVG PW=0.64U NW=0.42U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR4B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B2HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:38:10 2002                                       *
*******************************************************************************
.SUBCKT NOR4B2HD4X Z AN BN C D
MN4 Z NET17 GND GND N18 W=2.4U L=0.18U
MN3 Z NET47 GND GND N18 W=2.4U L=0.18U
MN2 Z D GND GND N18 W=2.4U L=0.18U
MN0 Z C GND GND N18 W=2.4U L=0.18U
MP4 NET37 D Z VDD P18 W=6.72U L=0.18U
MP3 NET27 C NET37 VDD P18 W=6.72U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=6.72U L=0.18U
MP2 NET12 NET47 NET27 VDD P18 W=6.72U L=0.18U
XI4 NET47 BN IVG PW=1.68U NW=1.12U
XI3 NET17 AN IVG PW=1.68U NW=1.12U
.ENDS NOR4B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B2HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:38:08 2002                                       *
*******************************************************************************
.SUBCKT NOR4B2HD2X Z AN BN C D
MN4 Z NET17 GND GND N18 W=1.2U L=0.18U
MN3 Z NET47 GND GND N18 W=1.2U L=0.18U
MN2 Z D GND GND N18 W=1.2U L=0.18U
MN0 Z C GND GND N18 W=1.2U L=0.18U
MP4 NET37 D Z VDD P18 W=3.36U L=0.18U
MP3 NET27 C NET37 VDD P18 W=3.36U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=3.36U L=0.18U
MP2 NET12 NET47 NET27 VDD P18 W=3.36U L=0.18U
XI4 NET47 BN IVG PW=1.12U NW=0.74U
XI3 NET17 AN IVG PW=1.12U NW=0.74U
.ENDS NOR4B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B2HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:38:06 2002                                       *
*******************************************************************************
.SUBCKT NOR4B2HD1X Z AN BN C D
MN4 Z NET17 GND GND N18 W=0.6U L=0.18U
MN3 Z NET47 GND GND N18 W=0.6U L=0.18U
MN2 Z D GND GND N18 W=0.6U L=0.18U
MN0 Z C GND GND N18 W=0.6U L=0.18U
MP4 NET37 D Z VDD P18 W=1.68U L=0.18U
MP3 NET27 C NET37 VDD P18 W=1.68U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 NET47 NET27 VDD P18 W=1.68U L=0.18U
XI4 NET47 BN IVG PW=0.64U NW=0.42U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR4B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B1HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:38:19 2002                                       *
*******************************************************************************
.SUBCKT NOR4B1HDLX Z AN B C D
MN4 Z NET17 GND GND N18 W=0.42U L=0.18U
MN3 Z B GND GND N18 W=0.42U L=0.18U
MN2 Z D GND GND N18 W=0.42U L=0.18U
MN0 Z C GND GND N18 W=0.42U L=0.18U
MP4 NET36 D Z VDD P18 W=1.16U L=0.18U
MP3 NET27 C NET36 VDD P18 W=1.16U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.16U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.16U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR4B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B1HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:38:18 2002                                       *
*******************************************************************************
.SUBCKT NOR4B1HD4X Z AN B C D
MN4 Z NET17 GND GND N18 W=2.4U L=0.18U
MN3 Z B GND GND N18 W=2.4U L=0.18U
MN2 Z D GND GND N18 W=2.4U L=0.18U
MN0 Z C GND GND N18 W=2.4U L=0.18U
MP4 NET36 D Z VDD P18 W=6.72U L=0.18U
MP3 NET27 C NET36 VDD P18 W=6.72U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=6.72U L=0.18U
MP2 NET12 B NET27 VDD P18 W=6.72U L=0.18U
XI3 NET17 AN IVG PW=1.68U NW=1.12U
.ENDS NOR4B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B1HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:38:16 2002                                       *
*******************************************************************************
.SUBCKT NOR4B1HD2X Z AN B C D
MN4 Z NET17 GND GND N18 W=1.2U L=0.18U
MN3 Z B GND GND N18 W=1.2U L=0.18U
MN2 Z D GND GND N18 W=1.2U L=0.18U
MN0 Z C GND GND N18 W=1.2U L=0.18U
MP4 NET36 D Z VDD P18 W=3.36U L=0.18U
MP3 NET27 C NET36 VDD P18 W=3.36U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=3.36U L=0.18U
MP2 NET12 B NET27 VDD P18 W=3.36U L=0.18U
XI3 NET17 AN IVG PW=1.12U NW=0.74U
.ENDS NOR4B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR4B1HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:38:14 2002                                       *
*******************************************************************************
.SUBCKT NOR4B1HD1X Z AN B C D
MN4 Z NET17 GND GND N18 W=0.6U L=0.18U
MN3 Z B GND GND N18 W=0.6U L=0.18U
MN2 Z D GND GND N18 W=0.6U L=0.18U
MN0 Z C GND GND N18 W=0.6U L=0.18U
MP4 NET36 D Z VDD P18 W=1.68U L=0.18U
MP3 NET27 C NET36 VDD P18 W=1.68U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR4B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:38:05 2002                                       *
*******************************************************************************
.SUBCKT NOR3HDLX Z A B C
MN3 Z A GND GND N18 W=0.42U L=0.18U
MN2 Z C GND GND N18 W=0.42U L=0.18U
MN0 Z B GND GND N18 W=0.42U L=0.18U
MP3 NET27 C Z VDD P18 W=1.0U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.0U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.0U L=0.18U
.ENDS NOR3HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:38:04 2002                                       *
*******************************************************************************
.SUBCKT NOR3HD4X Z A B C
MN3 Z A GND GND N18 W=2.8U L=0.18U
MN2 Z C GND GND N18 W=2.8U L=0.18U
MN0 Z B GND GND N18 W=2.8U L=0.18U
MP3 NET27 C Z VDD P18 W=6.72U L=0.18U
MP1 VDD A NET12 VDD P18 W=6.72U L=0.18U
MP2 NET12 B NET27 VDD P18 W=6.72U L=0.18U
.ENDS NOR3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:38:02 2002                                       *
*******************************************************************************
.SUBCKT NOR3HD2X Z A B C
MN3 Z A GND GND N18 W=1.4U L=0.18U
MN2 Z C GND GND N18 W=1.4U L=0.18U
MN0 Z B GND GND N18 W=1.4U L=0.18U
MP3 NET27 C Z VDD P18 W=3.36U L=0.18U
MP1 VDD A NET12 VDD P18 W=3.36U L=0.18U
MP2 NET12 B NET27 VDD P18 W=3.36U L=0.18U
.ENDS NOR3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:38:01 2002                                       *
*******************************************************************************
.SUBCKT NOR3HD1X Z A B C
MN3 Z A GND GND N18 W=0.7U L=0.18U
MN2 Z C GND GND N18 W=0.7U L=0.18U
MN0 Z B GND GND N18 W=0.7U L=0.18U
MP3 NET27 C Z VDD P18 W=1.68U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
.ENDS NOR3HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3B1HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:37:59 2002                                       *
*******************************************************************************
.SUBCKT NOR3B1HDLX Z AN B C
MN3 Z NET17 GND GND N18 W=0.42U L=0.18U
MN2 Z C GND GND N18 W=0.42U L=0.18U
MN0 Z B GND GND N18 W=0.42U L=0.18U
MP3 NET27 C Z VDD P18 W=1.0U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.0U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.0U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR3B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3B1HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:37:57 2002                                       *
*******************************************************************************
.SUBCKT NOR3B1HD4X Z AN B C
MN3 Z NET17 GND GND N18 W=2.8U L=0.18U
MN2 Z C GND GND N18 W=2.8U L=0.18U
MN0 Z B GND GND N18 W=2.8U L=0.18U
MP3 NET27 C Z VDD P18 W=6.72U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=6.72U L=0.18U
MP2 NET12 B NET27 VDD P18 W=6.72U L=0.18U
XI3 NET17 AN IVG PW=1.68U NW=1.12U
.ENDS NOR3B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3B1HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:37:55 2002                                       *
*******************************************************************************
.SUBCKT NOR3B1HD2X Z AN B C
MN3 Z NET17 GND GND N18 W=1.4U L=0.18U
MN2 Z C GND GND N18 W=1.4U L=0.18U
MN0 Z B GND GND N18 W=1.4U L=0.18U
MP3 NET27 C Z VDD P18 W=3.36U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=3.36U L=0.18U
MP2 NET12 B NET27 VDD P18 W=3.36U L=0.18U
XI3 NET17 AN IVG PW=1.12U NW=0.74U
.ENDS NOR3B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR3B1HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:37:54 2002                                       *
*******************************************************************************
.SUBCKT NOR3B1HD1X Z AN B C
MN3 Z NET17 GND GND N18 W=0.7U L=0.18U
MN2 Z C GND GND N18 W=0.7U L=0.18U
MN0 Z B GND GND N18 W=0.7U L=0.18U
MP3 NET27 C Z VDD P18 W=1.68U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.68U L=0.18U
MP2 NET12 B NET27 VDD P18 W=1.68U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR3B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:37:52 2002                                       *
*******************************************************************************
.SUBCKT NOR2HDLX Z A B
MN2 Z B GND GND N18 W=0.42U L=0.18U
MN0 Z A GND GND N18 W=0.42U L=0.18U
MP1 VDD A NET12 VDD P18 W=0.84U L=0.18U
MP2 NET12 B Z VDD P18 W=0.84U L=0.18U
.ENDS NOR2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HD4XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:37:51 2002                                       *
*******************************************************************************
.SUBCKT NOR2HD4XSPG Z A B
MN2 Z B GND GND N18 W=3.12U L=0.18U
MN0 Z A GND GND N18 W=3.12U L=0.18U
MP1 VDD A NET12 VDD P18 W=6.16U L=0.18U
MP2 NET12 B Z VDD P18 W=6.16U L=0.18U
.ENDS NOR2HD4XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:37:49 2002                                       *
*******************************************************************************
.SUBCKT NOR2HD4X Z A B
MN2 Z B GND GND N18 W=3.12U L=0.18U
MN0 Z A GND GND N18 W=3.12U L=0.18U
MP1 VDD A NET12 VDD P18 W=6.16U L=0.18U
MP2 NET12 B Z VDD P18 W=6.16U L=0.18U
.ENDS NOR2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HD2XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:37:47 2002                                       *
*******************************************************************************
.SUBCKT NOR2HD2XSPG Z A B
MN2 Z B GND GND N18 W=1.54U L=0.18U
MN0 Z A GND GND N18 W=1.54U L=0.18U
MP1 VDD A NET12 VDD P18 W=3.08U L=0.18U
MP2 NET12 B Z VDD P18 W=3.08U L=0.18U
.ENDS NOR2HD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:37:46 2002                                       *
*******************************************************************************
.SUBCKT NOR2HD2X Z A B
MN2 Z B GND GND N18 W=1.54U L=0.18U
MN0 Z A GND GND N18 W=1.54U L=0.18U
MP1 VDD A NET12 VDD P18 W=3.08U L=0.18U
MP2 NET12 B Z VDD P18 W=3.08U L=0.18U
.ENDS NOR2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:37:44 2002                                       *
*******************************************************************************
.SUBCKT NOR2HD1X Z A B
MN2 Z B GND GND N18 W=0.77U L=0.18U
MN0 Z A GND GND N18 W=0.77U L=0.18U
MP1 VDD A NET12 VDD P18 W=1.54U L=0.18U
MP2 NET12 B Z VDD P18 W=1.54U L=0.18U
.ENDS NOR2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2B1HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:37:42 2002                                       *
*******************************************************************************
.SUBCKT NOR2B1HDLX Z AN B
MN2 Z B GND GND N18 W=0.42U L=0.18U
MN0 Z NET17 GND GND N18 W=0.42U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=0.84U L=0.18U
MP2 NET12 B Z VDD P18 W=0.84U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR2B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2B1HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:37:40 2002                                       *
*******************************************************************************
.SUBCKT NOR2B1HD4X Z AN B
MN2 Z B GND GND N18 W=3.12U L=0.18U
MN0 Z NET17 GND GND N18 W=3.12U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=6.16U L=0.18U
MP2 NET12 B Z VDD P18 W=6.16U L=0.18U
XI3 NET17 AN IVG PW=1.68U NW=1.12U
.ENDS NOR2B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2B1HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:37:39 2002                                       *
*******************************************************************************
.SUBCKT NOR2B1HD2X Z AN B
MN2 Z B GND GND N18 W=1.54U L=0.18U
MN0 Z NET17 GND GND N18 W=1.54U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=3.08U L=0.18U
MP2 NET12 B Z VDD P18 W=3.08U L=0.18U
XI3 NET17 AN IVG PW=1.06U NW=0.7U
.ENDS NOR2B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NOR2B1HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:37:37 2002                                       *
*******************************************************************************
.SUBCKT NOR2B1HD1X Z AN B
MN2 Z B GND GND N18 W=0.77U L=0.18U
MN0 Z NET17 GND GND N18 W=0.77U L=0.18U
MP1 VDD NET17 NET12 VDD P18 W=1.54U L=0.18U
MP2 NET12 B Z VDD P18 W=1.54U L=0.18U
XI3 NET17 AN IVG PW=0.64U NW=0.42U
.ENDS NOR2B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:37:35 2002                                       *
*******************************************************************************
.SUBCKT NAND4HDLX Z A B C D
MN4 NET7 B NET25 GND N18 W=0.64U L=0.18U
MN5 NET25 A GND GND N18 W=0.64U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.64U L=0.18U
MN0 Z D NET10 GND N18 W=0.64U L=0.18U
MP3 VDD A Z VDD P18 W=0.64U L=0.18U
MP2 VDD D Z VDD P18 W=0.64U L=0.18U
MP1 VDD C Z VDD P18 W=0.64U L=0.18U
MP0 VDD B Z VDD P18 W=0.64U L=0.18U
.ENDS NAND4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:37:34 2002                                       *
*******************************************************************************
.SUBCKT NAND4HD4X Z A B C D
MN4 NET7 B NET25 GND N18 W=4.72U L=0.18U
MN5 NET25 A GND GND N18 W=4.72U L=0.18U
MN3 NET10 C NET7 GND N18 W=4.72U L=0.18U
MN0 Z D NET10 GND N18 W=4.72U L=0.18U
MP3 VDD A Z VDD P18 W=4.8U L=0.18U
MP2 VDD D Z VDD P18 W=4.8U L=0.18U
MP1 VDD C Z VDD P18 W=4.8U L=0.18U
MP0 VDD B Z VDD P18 W=4.8U L=0.18U
.ENDS NAND4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:37:32 2002                                       *
*******************************************************************************
.SUBCKT NAND4HD2X Z A B C D
MN4 NET7 B NET25 GND N18 W=2.36U L=0.18U
MN5 NET25 A GND GND N18 W=2.36U L=0.18U
MN3 NET10 C NET7 GND N18 W=2.36U L=0.18U
MN0 Z D NET10 GND N18 W=2.36U L=0.18U
MP3 VDD A Z VDD P18 W=2.4U L=0.18U
MP2 VDD D Z VDD P18 W=2.4U L=0.18U
MP1 VDD C Z VDD P18 W=2.4U L=0.18U
MP0 VDD B Z VDD P18 W=2.4U L=0.18U
.ENDS NAND4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:37:31 2002                                       *
*******************************************************************************
.SUBCKT NAND4HD1X Z A B C D
MN4 NET7 B NET25 GND N18 W=1.18U L=0.18U
MN5 NET25 A GND GND N18 W=1.18U L=0.18U
MN3 NET10 C NET7 GND N18 W=1.18U L=0.18U
MN0 Z D NET10 GND N18 W=1.18U L=0.18U
MP3 VDD A Z VDD P18 W=1.2U L=0.18U
MP2 VDD D Z VDD P18 W=1.2U L=0.18U
MP1 VDD C Z VDD P18 W=1.2U L=0.18U
MP0 VDD B Z VDD P18 W=1.2U L=0.18U
.ENDS NAND4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B2HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:37:23 2002                                       *
*******************************************************************************
.SUBCKT NAND4B2HDLX Z AN BN C D
XI5 NET39 BN IVG PW=0.64U NW=0.42U
XI4 NET42 AN IVG PW=0.64U NW=0.42U
MN4 NET7 NET39 NET32 GND N18 W=0.64U L=0.18U
MN5 NET32 NET42 GND GND N18 W=0.64U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.64U L=0.18U
MN0 Z D NET10 GND N18 W=0.64U L=0.18U
MP3 VDD NET42 Z VDD P18 W=0.64U L=0.18U
MP2 VDD D Z VDD P18 W=0.64U L=0.18U
MP1 VDD C Z VDD P18 W=0.64U L=0.18U
MP0 VDD NET39 Z VDD P18 W=0.64U L=0.18U
.ENDS NAND4B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B2HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:37:21 2002                                       *
*******************************************************************************
.SUBCKT NAND4B2HD4X Z AN BN C D
XI6 NET39 BN IVG PW=1.68U NW=1.12U
XI4 NET42 AN IVG PW=1.68U NW=1.12U
MN4 NET7 NET39 NET31 GND N18 W=4.72U L=0.18U
MN5 NET31 NET42 GND GND N18 W=4.72U L=0.18U
MN3 NET10 C NET7 GND N18 W=4.72U L=0.18U
MN0 Z D NET10 GND N18 W=4.72U L=0.18U
MP3 VDD NET42 Z VDD P18 W=4.8U L=0.18U
MP2 VDD D Z VDD P18 W=4.8U L=0.18U
MP1 VDD C Z VDD P18 W=4.8U L=0.18U
MP0 VDD NET39 Z VDD P18 W=4.8U L=0.18U
.ENDS NAND4B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B2HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:37:20 2002                                       *
*******************************************************************************
.SUBCKT NAND4B2HD2X Z AN BN C D
XI4 NET42 AN IVG PW=1.18U NW=0.78U
XI5 NET39 BN IVG PW=1.18U NW=0.78U
MN4 NET7 NET39 NET31 GND N18 W=2.36U L=0.18U
MN5 NET31 NET42 GND GND N18 W=2.36U L=0.18U
MN3 NET10 C NET7 GND N18 W=2.36U L=0.18U
MN0 Z D NET10 GND N18 W=2.36U L=0.18U
MP3 VDD NET42 Z VDD P18 W=2.4U L=0.18U
MP2 VDD D Z VDD P18 W=2.4U L=0.18U
MP1 VDD C Z VDD P18 W=2.4U L=0.18U
MP0 VDD NET39 Z VDD P18 W=2.4U L=0.18U
.ENDS NAND4B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B2HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:37:19 2002                                       *
*******************************************************************************
.SUBCKT NAND4B2HD1X Z AN BN C D
XI4 NET42 AN IVG PW=0.64U NW=0.42U
XI5 NET39 BN IVG PW=0.64U NW=0.42U
MN4 NET7 NET39 NET31 GND N18 W=1.18U L=0.18U
MN5 NET31 NET42 GND GND N18 W=1.18U L=0.18U
MN3 NET10 C NET7 GND N18 W=1.18U L=0.18U
MN0 Z D NET10 GND N18 W=1.18U L=0.18U
MP3 VDD NET42 Z VDD P18 W=1.2U L=0.18U
MP2 VDD D Z VDD P18 W=1.2U L=0.18U
MP1 VDD C Z VDD P18 W=1.2U L=0.18U
MP0 VDD NET39 Z VDD P18 W=1.2U L=0.18U
.ENDS NAND4B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B1HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:37:28 2002                                       *
*******************************************************************************
.SUBCKT NAND4B1HDLX Z AN B C D
XI3 NET36 AN IVG PW=0.64U NW=0.42U
MN4 NET7 B NET28 GND N18 W=0.64U L=0.18U
MN5 NET28 NET36 GND GND N18 W=0.64U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.64U L=0.18U
MN0 Z D NET10 GND N18 W=0.64U L=0.18U
MP3 VDD NET36 Z VDD P18 W=0.64U L=0.18U
MP2 VDD D Z VDD P18 W=0.64U L=0.18U
MP1 VDD C Z VDD P18 W=0.64U L=0.18U
MP0 VDD B Z VDD P18 W=0.64U L=0.18U
.ENDS NAND4B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B1HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:37:28 2002                                       *
*******************************************************************************
.SUBCKT NAND4B1HD4X Z AN B C D
XI3 NET36 AN IVG PW=1.68U NW=1.12U
MN4 NET7 B NET28 GND N18 W=4.72U L=0.18U
MN5 NET28 NET36 GND GND N18 W=4.72U L=0.18U
MN3 NET10 C NET7 GND N18 W=4.72U L=0.18U
MN0 Z D NET10 GND N18 W=4.72U L=0.18U
MP3 VDD NET36 Z VDD P18 W=4.8U L=0.18U
MP2 VDD D Z VDD P18 W=4.8U L=0.18U
MP1 VDD C Z VDD P18 W=4.8U L=0.18U
MP0 VDD B Z VDD P18 W=4.8U L=0.18U
.ENDS NAND4B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B1HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:37:25 2002                                       *
*******************************************************************************
.SUBCKT NAND4B1HD2X Z AN B C D
XI3 NET36 AN IVG PW=1.18U NW=0.78U
MN4 NET7 B NET28 GND N18 W=2.36U L=0.18U
MN5 NET28 NET36 GND GND N18 W=2.36U L=0.18U
MN3 NET10 C NET7 GND N18 W=2.36U L=0.18U
MN0 Z D NET10 GND N18 W=2.36U L=0.18U
MP3 VDD NET36 Z VDD P18 W=2.4U L=0.18U
MP2 VDD D Z VDD P18 W=2.4U L=0.18U
MP1 VDD C Z VDD P18 W=2.4U L=0.18U
MP0 VDD B Z VDD P18 W=2.4U L=0.18U
.ENDS NAND4B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND4B1HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:37:24 2002                                       *
*******************************************************************************
.SUBCKT NAND4B1HD1X Z AN B C D
XI3 NET36 AN IVG PW=0.64U NW=0.42U
MN4 NET7 B NET28 GND N18 W=1.18U L=0.18U
MN5 NET28 NET36 GND GND N18 W=1.18U L=0.18U
MN3 NET10 C NET7 GND N18 W=1.18U L=0.18U
MN0 Z D NET10 GND N18 W=1.18U L=0.18U
MP3 VDD NET36 Z VDD P18 W=1.2U L=0.18U
MP2 VDD D Z VDD P18 W=1.2U L=0.18U
MP1 VDD C Z VDD P18 W=1.2U L=0.18U
MP0 VDD B Z VDD P18 W=1.2U L=0.18U
.ENDS NAND4B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3ODHD                                                            *
* LAST TIME SAVED: AUG 30 10:37:09 2002                                       *
*******************************************************************************
.SUBCKT NAND3ODHD Z A B C
MP4 VDD C NET9 VDD P18 W=0.64U L=0.18U
MP3 VDD NET9 NET22 VDD P18 W=1.68U L=0.18U
MP0 VDD A NET9 VDD P18 W=0.64U L=0.18U
MP1 VDD B NET9 VDD P18 W=0.64U L=0.18U
MN5 NET9 C NET43 GND N18 W=0.58U L=0.18U
MN2 Z NET22 GND GND N18 W=1.18U L=0.18U M=2
MN1 NET22 NET9 GND GND N18 W=0.84U L=0.18U
MN3 NET43 B NET31 GND N18 W=0.58U L=0.18U
MN4 NET31 A GND GND N18 W=0.58U L=0.18U
.ENDS NAND3ODHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:37:17 2002                                       *
*******************************************************************************
.SUBCKT NAND3HDLX Z A B C
MN4 NET7 A GND GND N18 W=0.58U L=0.18U
MN3 NET10 B NET7 GND N18 W=0.58U L=0.18U
MN0 Z C NET10 GND N18 W=0.58U L=0.18U
MP2 VDD C Z VDD P18 W=0.64U L=0.18U
MP1 VDD B Z VDD P18 W=0.64U L=0.18U
MP0 VDD A Z VDD P18 W=0.64U L=0.18U
.ENDS NAND3HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:37:15 2002                                       *
*******************************************************************************
.SUBCKT NAND3HD4X Z A B C
MN4 NET7 A GND GND N18 W=4.4U L=0.18U
MN3 NET10 B NET7 GND N18 W=4.4U L=0.18U
MN0 Z C NET10 GND N18 W=4.4U L=0.18U
MP2 VDD C Z VDD P18 W=4.8U L=0.18U
MP1 VDD B Z VDD P18 W=4.8U L=0.18U
MP0 VDD A Z VDD P18 W=4.8U L=0.18U
.ENDS NAND3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:37:14 2002                                       *
*******************************************************************************
.SUBCKT NAND3HD2X Z A B C
MN4 NET7 A GND GND N18 W=2.2U L=0.18U
MN3 NET10 B NET7 GND N18 W=2.2U L=0.18U
MN0 Z C NET10 GND N18 W=2.2U L=0.18U
MP2 VDD C Z VDD P18 W=2.4U L=0.18U
MP1 VDD B Z VDD P18 W=2.4U L=0.18U
MP0 VDD A Z VDD P18 W=2.4U L=0.18U
.ENDS NAND3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:37:12 2002                                       *
*******************************************************************************
.SUBCKT NAND3HD1X Z A B C
MN4 NET7 A GND GND N18 W=1.1U L=0.18U
MN3 NET10 B NET7 GND N18 W=1.1U L=0.18U
MN0 Z C NET10 GND N18 W=1.1U L=0.18U
MP2 VDD C Z VDD P18 W=1.2U L=0.18U
MP1 VDD B Z VDD P18 W=1.2U L=0.18U
MP0 VDD A Z VDD P18 W=1.2U L=0.18U
.ENDS NAND3HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3B1HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:37:09 2002                                       *
*******************************************************************************
.SUBCKT NAND3B1HDLX Z AN B C
XI3 NET20 AN IVG PW=0.64U NW=0.42U
MN4 NET7 NET20 GND GND N18 W=0.58U L=0.18U
MN3 NET10 B NET7 GND N18 W=0.58U L=0.18U
MN0 Z C NET10 GND N18 W=0.58U L=0.18U
MP2 VDD C Z VDD P18 W=0.64U L=0.18U
MP1 VDD B Z VDD P18 W=0.64U L=0.18U
MP0 VDD NET20 Z VDD P18 W=0.64U L=0.18U
.ENDS NAND3B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3B1HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:37:07 2002                                       *
*******************************************************************************
.SUBCKT NAND3B1HD4X Z AN B C
XI3 NET20 AN IVG PW=1.68U NW=1.12U
MN4 NET7 NET20 GND GND N18 W=4.4U L=0.18U
MN3 NET10 B NET7 GND N18 W=4.4U L=0.18U
MN0 Z C NET10 GND N18 W=4.4U L=0.18U
MP2 VDD C Z VDD P18 W=4.8U L=0.18U
MP1 VDD B Z VDD P18 W=4.8U L=0.18U
MP0 VDD NET20 Z VDD P18 W=4.8U L=0.18U
.ENDS NAND3B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3B1HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:37:05 2002                                       *
*******************************************************************************
.SUBCKT NAND3B1HD2X Z AN B C
XI3 NET20 AN IVG PW=1.11U NW=0.74U
MN4 NET7 NET20 GND GND N18 W=2.2U L=0.18U
MN3 NET10 B NET7 GND N18 W=2.2U L=0.18U
MN0 Z C NET10 GND N18 W=2.2U L=0.18U
MP2 VDD C Z VDD P18 W=2.4U L=0.18U
MP1 VDD B Z VDD P18 W=2.4U L=0.18U
MP0 VDD NET20 Z VDD P18 W=2.4U L=0.18U
.ENDS NAND3B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND3B1HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:37:04 2002                                       *
*******************************************************************************
.SUBCKT NAND3B1HD1X Z AN B C
XI3 NET20 AN IVG PW=0.64U NW=0.42U
MN4 NET7 NET20 GND GND N18 W=1.1U L=0.18U
MN3 NET10 B NET7 GND N18 W=1.1U L=0.18U
MN0 Z C NET10 GND N18 W=1.1U L=0.18U
MP2 VDD C Z VDD P18 W=1.2U L=0.18U
MP1 VDD B Z VDD P18 W=1.2U L=0.18U
MP0 VDD NET20 Z VDD P18 W=1.2U L=0.18U
.ENDS NAND3B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2ODHD                                                            *
* LAST TIME SAVED: AUG 30 10:36:52 2002                                       *
*******************************************************************************
.SUBCKT NAND2ODHD Z A B
MP3 VDD NET9 NET22 VDD P18 W=1.68U L=0.18U
MP0 VDD A NET9 VDD P18 W=0.64U L=0.18U
MP1 VDD B NET9 VDD P18 W=0.64U L=0.18U
MN2 Z NET22 GND GND N18 W=1.18U L=0.18U M=2
MN1 NET22 NET9 GND GND N18 W=0.84U L=0.18U
MN3 NET9 B NET31 GND N18 W=0.52U L=0.18U
MN4 NET31 A GND GND N18 W=0.52U L=0.18U
.ENDS NAND2ODHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:37:02 2002                                       *
*******************************************************************************
.SUBCKT NAND2HDLX Z A B
MN1 NET6 A GND GND N18 W=0.54U L=0.18U
MN0 Z B NET6 GND N18 W=0.54U L=0.18U
MP1 VDD B Z VDD P18 W=0.64U L=0.18U
MP0 VDD A Z VDD P18 W=0.64U L=0.18U
.ENDS NAND2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HD4XSPG                                                         *
* LAST TIME SAVED: AUG 30 10:37:01 2002                                       *
*******************************************************************************
.SUBCKT NAND2HD4XSPG Z A B
MN1 NET6 A GND GND N18 W=3.66U L=0.18U
MN0 Z B NET6 GND N18 W=3.66U L=0.18U
MP1 VDD B Z VDD P18 W=4.8U L=0.18U
MP0 VDD A Z VDD P18 W=4.8U L=0.18U
.ENDS NAND2HD4XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:36:59 2002                                       *
*******************************************************************************
.SUBCKT NAND2HD4X Z A B
MN1 NET6 A GND GND N18 W=3.66U L=0.18U
MN0 Z B NET6 GND N18 W=3.66U L=0.18U
MP1 VDD B Z VDD P18 W=4.8U L=0.18U
MP0 VDD A Z VDD P18 W=4.8U L=0.18U
.ENDS NAND2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HD2XSPG                                                         *
* LAST TIME SAVED: AUG 30 10:36:57 2002                                       *
*******************************************************************************
.SUBCKT NAND2HD2XSPG Z A B
MN1 NET6 A GND GND N18 W=2.0U L=0.18U
MN0 Z B NET6 GND N18 W=2.0U L=0.18U
MP1 VDD B Z VDD P18 W=2.4U L=0.18U
MP0 VDD A Z VDD P18 W=2.4U L=0.18U
.ENDS NAND2HD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:36:56 2002                                       *
*******************************************************************************
.SUBCKT NAND2HD2X Z A B
MN1 NET6 A GND GND N18 W=2.0U L=0.18U
MN0 Z B NET6 GND N18 W=2.0U L=0.18U
MP1 VDD B Z VDD P18 W=2.4U L=0.18U
MP0 VDD A Z VDD P18 W=2.4U L=0.18U
.ENDS NAND2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:36:54 2002                                       *
*******************************************************************************
.SUBCKT NAND2HD1X Z A B
MN1 NET6 A GND GND N18 W=1.0U L=0.18U
MN0 Z B NET6 GND N18 W=1.0U L=0.18U
MP1 VDD B Z VDD P18 W=1.2U L=0.18U
MP0 VDD A Z VDD P18 W=1.2U L=0.18U
.ENDS NAND2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2B1HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:36:51 2002                                       *
*******************************************************************************
.SUBCKT NAND2B1HDLX Z AN B
XI3 NET14 AN IVG PW=0.64U NW=0.42U
MN1 NET6 NET14 GND GND N18 W=0.54U L=0.18U
MN0 Z B NET6 GND N18 W=0.54U L=0.18U
MP1 VDD NET14 Z VDD P18 W=0.64U L=0.18U
MP0 VDD B Z VDD P18 W=0.64U L=0.18U
.ENDS NAND2B1HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2B1HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:36:49 2002                                       *
*******************************************************************************
.SUBCKT NAND2B1HD4X Z AN B
XI3 NET14 AN IVG PW=1.68U NW=1.12U
MN1 NET6 NET14 GND GND N18 W=3.66U L=0.18U
MN0 Z B NET6 GND N18 W=3.66U L=0.18U
MP1 VDD NET14 Z VDD P18 W=4.8U L=0.18U
MP0 VDD B Z VDD P18 W=4.8U L=0.18U
.ENDS NAND2B1HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2B1HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:36:47 2002                                       *
*******************************************************************************
.SUBCKT NAND2B1HD2X Z AN B
XI3 NET14 AN IVG PW=1.0U NW=0.66U
MN1 NET6 NET14 GND GND N18 W=2.0U L=0.18U
MN0 Z B NET6 GND N18 W=2.0U L=0.18U
MP1 VDD NET14 Z VDD P18 W=2.4U L=0.18U
MP0 VDD B Z VDD P18 W=2.4U L=0.18U
.ENDS NAND2B1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: NAND2B1HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:36:45 2002                                       *
*******************************************************************************
.SUBCKT NAND2B1HD1X Z AN B
XI4 NET14 AN IVG PW=0.64U NW=0.42U
MN1 NET6 NET14 GND GND N18 W=1.0U L=0.18U
MN0 Z B NET6 GND N18 W=1.0U L=0.18U
MP1 VDD NET14 Z VDD P18 W=1.2U L=0.18U
MP0 VDD B Z VDD P18 W=1.2U L=0.18U
.ENDS NAND2B1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI4HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:36:43 2002                                       *
*******************************************************************************
.SUBCKT MUXI4HDLX Z A B C D S0 S1
XI7 NET39 NET14 NET45 S0 TG1G NW=0.42U PW=0.42U
XI10 NET33 NET26 S0 NET45 TG1G NW=0.42U PW=0.42U
XI4 NET49 NET18 S1 NET37 TG1G NW=0.42U PW=0.42U
XI11 NET47 NET18 NET37 S1 TG1G NW=0.42U PW=0.42U
XI5 NET43 NET14 S0 NET45 TG1G NW=0.42U PW=0.42U
XI9 NET35 NET26 NET45 S0 TG1G NW=0.42U PW=0.42U
XI12 NET37 S1 IVG PW=0.45U NW=0.3U
XI2 NET35 C IVG PW=0.45U NW=0.3U
XI8 NET39 A IVG PW=0.45U NW=0.3U
XI6 Z NET18 IVG PW=0.64U NW=0.42U
XI3 NET33 D IVG PW=0.45U NW=0.3U
XI1 NET43 B IVG PW=0.45U NW=0.3U
XI0 NET45 S0 IVG PW=0.64U NW=0.42U
XI16 NET47 NET14 IVG PW=0.64U NW=0.42U
XI17 NET49 NET26 IVG PW=0.64U NW=0.42U
.ENDS MUXI4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI4HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:36:41 2002                                       *
*******************************************************************************
.SUBCKT MUXI4HD4X Z A B C D S0 S1
XI16 NET15 NET36 IVG PW=1.68U NW=1.18U
XI6 Z NET48 IVG PW=4.8U NW=3.2U
XI12 NET19 S1 IVG PW=0.64U NW=0.42U
XI0 NET21 S0 IVG PW=1.14U NW=0.76U
XI8 NET23 A IVG PW=1.72U NW=1.2U
XI3 NET9 D IVG PW=1.72U NW=1.2U
XI2 NET11 C IVG PW=1.72U NW=1.2U
XI1 NET13 B IVG PW=1.72U NW=1.2U
XI13 NET25 NET44 IVG PW=1.68U NW=1.18U
XI11 NET15 NET48 NET19 S1 TG1G NW=1.18U PW=1.2U
XI7 NET23 NET36 NET21 S0 TG1G NW=1.0U PW=1.0U
XI14 NET13 NET36 S0 NET21 TG1G NW=1.0U PW=1.0U
XI15 NET11 NET44 NET21 S0 TG1G NW=1.0U PW=1.0U
XI17 NET9 NET44 S0 NET21 TG1G NW=1.0U PW=1.0U
XI18 NET25 NET48 S1 NET19 TG1G NW=1.18U PW=1.2U
.ENDS MUXI4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI4HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:36:39 2002                                       *
*******************************************************************************
.SUBCKT MUXI4HD2X Z A B C D S0 S1
XI7 NET41 NET22 NET43 S0 TG1G NW=1.0U PW=1.0U
XI14 NET39 NET22 S0 NET43 TG1G NW=1.0U PW=1.0U
XI15 NET37 NET14 NET43 S0 TG1G NW=1.0U PW=1.0U
XI17 NET35 NET14 S0 NET43 TG1G NW=1.0U PW=1.0U
XI18 NET33 NET10 S1 NET45 TG1G NW=1.18U PW=1.2U
XI20 NET49 NET10 NET45 S1 TG1G NW=1.18U PW=1.2U
XI8 NET41 A IVG PW=1.44U NW=0.97U
XI0 NET43 S0 IVG PW=0.9U NW=0.6U
XI3 NET35 D IVG PW=1.44U NW=0.97U
XI2 NET37 C IVG PW=1.44U NW=0.97U
XI1 NET39 B IVG PW=1.44U NW=0.97U
XI12 NET45 S1 IVG PW=0.64U NW=0.42U
XI6 Z NET10 IVG PW=2.4U NW=1.6U
XI16 NET49 NET22 IVG PW=1.68U NW=1.22U
XI19 NET33 NET14 IVG PW=1.68U NW=1.22U
.ENDS MUXI4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI4HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:36:37 2002                                       *
*******************************************************************************
.SUBCKT MUXI4HD1X Z A B C D S0 S1
XI17 NET9 NET36 IVG PW=0.9U NW=0.6U
XI16 NET11 NET44 IVG PW=0.9U NW=0.6U
XI0 NET23 S0 IVG PW=0.88U NW=0.58U
XI1 NET21 B IVG PW=0.72U NW=0.48U
XI2 NET19 C IVG PW=0.72U NW=0.48U
XI6 Z NET32 IVG PW=1.2U NW=0.8U
XI8 NET25 A IVG PW=0.72U NW=0.48U
XI9 NET17 D IVG PW=0.72U NW=0.48U
XI12 NET15 S1 IVG PW=0.45U NW=0.3U
XI14 NET19 NET36 NET23 S0 TG1G NW=0.6U PW=0.6U
XI15 NET17 NET36 S0 NET23 TG1G NW=0.6U PW=0.6U
XI11 NET11 NET32 NET15 S1 TG1G NW=0.6U PW=0.6U
XI10 NET9 NET32 S1 NET15 TG1G NW=0.6U PW=0.6U
XI13 NET21 NET44 S0 NET23 TG1G NW=0.6U PW=0.6U
XI7 NET25 NET44 NET23 S0 TG1G NW=0.6U PW=0.6U
.ENDS MUXI4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI2HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:36:35 2002                                       *
*******************************************************************************
.SUBCKT MUXI2HDLX Z A B S0
XI1 Z NET28 IVG PW=0.64U NW=0.42U
XI0 NET6 S0 IVG PW=0.45U NW=0.3U
XI4 A NET28 NET6 S0 TG1G NW=0.42U PW=0.42U
XI2 B NET28 S0 NET6 TG1G NW=0.42U PW=0.42U
.ENDS MUXI2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI2HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:36:34 2002                                       *
*******************************************************************************
.SUBCKT MUXI2HD4X Z A B S0
XI1 Z NET28 IVG PW=4.8U NW=3.2U
XI0 NET6 S0 IVG PW=0.64U NW=0.42U
XI4 A NET28 NET6 S0 TG1G NW=1.18U PW=1.2U
XI2 B NET28 S0 NET6 TG1G NW=1.18U PW=1.2U
.ENDS MUXI2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI2HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:36:32 2002                                       *
*******************************************************************************
.SUBCKT MUXI2HD2X Z A B S0
XI1 Z NET27 IVG PW=2.4U NW=1.6U
XI0 NET6 S0 IVG PW=0.64U NW=0.42U
XI4 A NET27 NET6 S0 TG1G NW=1.18U PW=1.2U
XI2 B NET27 S0 NET6 TG1G NW=1.18U PW=1.2U
.ENDS MUXI2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUXI2HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:36:30 2002                                       *
*******************************************************************************
.SUBCKT MUXI2HD1X Z A B S0
XI5 B NET13 S0 NET20 TG1G NW=0.6U PW=0.6U
XI4 A NET13 NET20 S0 TG1G NW=0.6U PW=0.6U
XI1 Z NET13 IVG PW=1.2U NW=0.8U
XI0 NET20 S0 IVG PW=0.45U NW=0.3U
.ENDS MUXI2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX4HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:36:29 2002                                       *
*******************************************************************************
.SUBCKT MUX4HDLX Z A B C D S0 S1
XI0 NET9 S0 IVG PW=0.64U NW=0.42U
XI13 NET17 B IVG PW=0.64U NW=0.42U
XI14 NET13 C IVG PW=0.64U NW=0.42U
XI8 NET15 A IVG PW=0.64U NW=0.42U
XI15 NET11 D IVG PW=0.64U NW=0.42U
XI6 Z NET40 IVG PW=0.64U NW=0.42U
XI12 NET21 S1 IVG PW=0.45U NW=0.3U
XI10 NET32 NET40 NET21 S1 TG1G NW=0.6U PW=0.6U
XI5 NET11 NET28 S0 NET9 TG1G NW=0.6U PW=0.6U
XI11 NET28 NET40 S1 NET21 TG1G NW=0.6U PW=0.6U
XI7 NET15 NET32 NET9 S0 TG1G NW=0.6U PW=0.6U
XI4 NET13 NET28 NET9 S0 TG1G NW=0.6U PW=0.6U
XI3 NET17 NET32 S0 NET9 TG1G NW=0.6U PW=0.6U
.ENDS MUX4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX4HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:36:27 2002                                       *
*******************************************************************************
.SUBCKT MUX4HD4X Z A B C D S0 S1
XI3 NET79 NET62 S0 NET81 TG1G NW=1.22U PW=1.72U
XI4 NET77 NET50 NET81 S0 TG1G NW=1.22U PW=1.72U
XI7 NET75 NET62 NET81 S0 TG1G NW=1.22U PW=1.72U
XI5 NET73 NET50 S0 NET81 TG1G NW=1.22U PW=1.72U
XI10 NET62 NET66 NET69 S1 TG1G NW=1.22U PW=1.72U
XI11 NET50 NET66 S1 NET69 TG1G NW=1.22U PW=1.72U
XI14 NET77 C IVG PW=1.72U NW=1.22U
XI0 NET81 S0 IVG PW=1.44U NW=0.96U
XI8 NET75 A IVG PW=1.72U NW=1.22U
XI15 NET73 D IVG PW=1.72U NW=1.22U
XI6 Z NET66 IVG PW=4.8U NW=3.2U
XI12 NET69 S1 IVG PW=0.72U NW=0.48U
XI13 NET79 B IVG PW=1.72U NW=1.22U
.ENDS MUX4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX4HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:36:25 2002                                       *
*******************************************************************************
.SUBCKT MUX4HD2X Z A B C D S0 S1
XI0 NET9 S0 IVG PW=1.44U NW=0.96U
XI13 NET17 B IVG PW=1.72U NW=1.22U
XI14 NET13 C IVG PW=1.72U NW=1.22U
XI8 NET15 A IVG PW=1.72U NW=1.22U
XI15 NET11 D IVG PW=1.72U NW=1.22U
XI6 Z NET40 IVG PW=2.4U NW=1.6U
XI12 NET21 S1 IVG PW=0.72U NW=0.48U
XI11 NET28 NET40 S1 NET21 TG1G NW=1.22U PW=1.72U
XI3 NET17 NET32 S0 NET9 TG1G NW=1.22U PW=1.72U
XI4 NET13 NET28 NET9 S0 TG1G NW=1.22U PW=1.72U
XI7 NET15 NET32 NET9 S0 TG1G NW=1.22U PW=1.72U
XI5 NET11 NET28 S0 NET9 TG1G NW=1.22U PW=1.72U
XI10 NET32 NET40 NET21 S1 TG1G NW=1.22U PW=1.72U
.ENDS MUX4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX4HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:36:23 2002                                       *
*******************************************************************************
.SUBCKT MUX4HD1X Z A B C D S0 S1
XI7 NET26 NET9 NET34 S0 TG1G NW=1.18U PW=1.2U
XI22 NET28 NET82 NET34 S0 TG1G NW=1.18U PW=1.2U
XI25 NET82 NET17 S1 NET89 TG1G NW=1.18U PW=1.2U
XI24 NET9 NET17 NET89 S1 TG1G NW=1.18U PW=1.2U
XI23 NET32 NET82 S0 NET34 TG1G NW=1.18U PW=1.2U
XI21 NET24 NET9 S0 NET34 TG1G NW=1.18U PW=1.2U
XI12 NET89 S1 IVG PW=0.64U NW=0.42U
XI20 NET32 D IVG PW=1.44U NW=0.97U
XI8 NET26 A IVG PW=1.44U NW=0.97U
XI6 Z NET17 IVG PW=1.2U NW=0.8U
XI19 NET28 C IVG PW=1.44U NW=0.97U
XI18 NET24 B IVG PW=1.44U NW=0.97U
XI0 NET34 S0 IVG PW=0.88U NW=0.58U
.ENDS MUX4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX2HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:36:22 2002                                       *
*******************************************************************************
.SUBCKT MUX2HDLX Z A B S0
XI5 NET18 NET7 S0 NET20 TG1G NW=0.42U PW=0.42U
XI4 NET16 NET7 NET20 S0 TG1G NW=0.42U PW=0.42U
XI6 Z NET7 IVG PW=0.64U NW=0.42U
XI3 NET16 A IVG PW=0.64U NW=0.42U
XI2 NET18 B IVG PW=0.64U NW=0.42U
XI0 NET20 S0 IVG PW=0.45U NW=0.3U
.ENDS MUX2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX2HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:36:20 2002                                       *
*******************************************************************************
.SUBCKT MUX2HD4X Z A B S0
XI9 Z NET15 IVG PW=4.8U NW=3.2U
XI8 NET8 A IVG PW=1.68U NW=1.18U
XI12 NET10 B IVG PW=1.68U NW=1.18U
XI13 NET12 S0 IVG PW=0.64U NW=0.42U
XI11 NET10 NET15 S0 NET12 TG1G NW=1.18U PW=1.2U
XI10 NET8 NET15 NET12 S0 TG1G NW=1.18U PW=1.2U
.ENDS MUX2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX2HD2XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:36:18 2002                                       *
*******************************************************************************
.SUBCKT MUX2HD2XSPG Z A B S0
XI7 NET18 NET11 NET14 S0 TG1G NW=1.18U PW=1.2U
XI13 NET16 NET11 S0 NET14 TG1G NW=1.18U PW=1.2U
XI11 NET14 S0 IVG PW=0.64U NW=0.42U
XI9 NET18 A IVG PW=1.68U NW=1.18U
XI8 Z NET11 IVG PW=2.4U NW=1.6U
XI12 NET16 B IVG PW=1.68U NW=1.18U
.ENDS MUX2HD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX2HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:36:17 2002                                       *
*******************************************************************************
.SUBCKT MUX2HD2X Z A B S0
XI7 NET18 NET11 NET14 S0 TG1G NW=1.18U PW=1.2U
XI13 NET16 NET11 S0 NET14 TG1G NW=1.18U PW=1.2U
XI11 NET14 S0 IVG PW=0.64U NW=0.42U
XI9 NET18 A IVG PW=1.68U NW=1.18U
XI8 Z NET11 IVG PW=2.4U NW=1.6U
XI12 NET16 B IVG PW=1.68U NW=1.18U
.ENDS MUX2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MUX2HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:36:15 2002                                       *
*******************************************************************************
.SUBCKT MUX2HD1X Z A B S0
XI0 NET6 S0 IVG PW=0.45U NW=0.3U
XI1 NET8 B IVG PW=0.9U NW=0.6U
XI3 NET10 A IVG PW=0.9U NW=0.6U
XI6 Z NET19 IVG PW=1.2U NW=0.8U
XI4 NET10 NET19 NET6 S0 TG1G NW=0.6U PW=0.6U
XI5 NET8 NET19 S0 NET6 TG1G NW=0.6U PW=0.6U
.ENDS MUX2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRIIVG                                                               *
* LAST TIME SAVED: SEP 12 11:15:39 2001                                       *
*******************************************************************************
.SUBCKT TRIIVG Z A CK CKN NL=0.18U NW=0.24U PL=0.18U PW=0.24U
MP1 VDD A NET16 VDD P18 W=PW L=PL
MP0 NET16 CKN Z VDD P18 W=PW L=PL
MN0 Z CK NET18 GND N18 W=NW L=NL
MN1 GND A NET18 GND N18 W=NW L=NL
.ENDS TRIIVG

*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRIIVG_1                                                             *
* LAST TIME SAVED: SEP 12 11:15:39 2001                                       *
*******************************************************************************
.SUBCKT TRIIVG_1 Z A CK CKN NL0=0.18U NL1=0.18U NW=0.24U PL0=0.18U PL1=0.18U PW=0.24U
MP1 VDD A NET16 VDD P18 W=PW L=PL1
MP0 NET16 CKN Z VDD P18 W=PW L=PL0
MN0 Z CK NET18 GND N18 W=NW L=NL0
MN1 GND A NET18 GND N18 W=NW L=NL1
.ENDS TRIIVG_1



*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATTSHDLX                                                            *
* LAST TIME SAVED: MAR  4 16:21:28 2003                                       *
*******************************************************************************
.SUBCKT LATTSHDLX Q D E G
XI11 NET31 NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI20 Q NETQ E NET20 TRIIVG NW=0.8U PW=1.2U
XI9 D NET31 NET24 NET32 TG1G NW=0.7U PW=0.7U
XI19 NET20 E IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI10 NETQ NET31 IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATTSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD4X                                                            *
* LAST TIME SAVED: AUG 30 10:44:34 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD4X Z A E
MN0 Z NET9 GND GND N18 W=3.2U L=0.18U
MN1 NET9 A GND GND N18 W=1.2U L=0.18U
MN2 NET9 NET27 GND GND N18 W=0.42U L=0.18U
MP0 VDD A NET14 VDD P18 W=1.72U L=0.18U
MP1 VDD E NET14 VDD P18 W=0.64U L=0.18U
MP4 VDD NET14 Z VDD P18 W=4.8U L=0.18U
XI6 NET9 NET14 E NET27 TG1G NW=0.7U PW=0.7U
XI3 NET27 E IVG PW=0.45U NW=0.30U
.ENDS BUFTSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATTSHD4X                                                            *
* LAST TIME SAVED: MAR  4 16:21:12 2003                                       *
*******************************************************************************
.SUBCKT LATTSHD4X Q D E G
XI23 Q NETQ E BUFTSHD4X
XI11 NETQ NET27 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI10 NET27 NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATTSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD2X                                                            *
* LAST TIME SAVED: AUG 30 10:44:15 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD2X Z A E
MN1 NET9 A GND GND N18 W=0.56U L=0.18U
MN2 NET9 NET27 GND GND N18 W=0.42U L=0.18U
MN0 Z NET9 GND GND N18 W=1.6U L=0.18U
MP1 VDD E NET14 VDD P18 W=0.6U L=0.18U
MP4 VDD NET14 Z VDD P18 W=2.4U L=0.18U
MP0 VDD A NET14 VDD P18 W=0.96U L=0.18U
XI6 NET9 NET14 E NET27 TG1G NW=0.4U PW=0.4U
XI3 NET27 E IVG PW=0.45U NW=0.30U
.ENDS BUFTSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATTSHD2X                                                            *
* LAST TIME SAVED: MAR  4 16:20:56 2003                                       *
*******************************************************************************
.SUBCKT LATTSHD2X Q D E G
XI23 Q NETQ E BUFTSHD2X
XI11 NETQ NET27 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI10 NET27 NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATTSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATTSHD1X                                                            *
* LAST TIME SAVED: MAR  4 16:20:41 2003                                       *
*******************************************************************************
.SUBCKT LATTSHD1X Q D E G
XI11 NET31 NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI20 Q NETQ E NET20 TRIIVG NW=1.22U PW=1.72U
XI9 D NET31 NET24 NET32 TG1G NW=0.7U PW=0.7U
XI19 NET20 E IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI10 NETQ NET31 IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATTSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSRHDLX                                                            *
* LAST TIME SAVED: MAR  4 16:20:27 2003                                       *
*******************************************************************************
.SUBCKT LATSRHDLX Q QN D G RN SN
MP8 VDD RN NET52 VDD P18 W=0.84U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.16U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.16U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NETQ VDD P18 W=0.84U L=0.18U
MN6 NETQ NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=0.77U L=0.18U
MN2 NET47 D NET44 GND N18 W=0.77U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET80 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSRHD4X                                                            *
* LAST TIME SAVED: MAR  4 16:20:11 2003                                       *
*******************************************************************************
.SUBCKT LATSRHD4X Q QN D G RN SN
MP8 VDD RN NET52 VDD P18 W=1.44U L=0.18U
MP6 NET103 D NET47 VDD P18 W=3.3U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=3.3U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1.68U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NETQ VDD P18 W=1.44U L=0.18U
MN6 NETQ NET80 GND GND N18 W=0.72U L=0.18U
MN3 NET44 RN GND GND N18 W=2.3U L=0.18U
MN2 NET47 D NET44 GND N18 W=2.3U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.8U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=1.18U PW=1.18U
XI21 NET80 SN IVG PW=1.5U NW=1U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSRHD2X                                                            *
* LAST TIME SAVED: MAR  4 16:19:27 2003                                       *
*******************************************************************************
.SUBCKT LATSRHD2X Q QN D G RN SN
MP8 VDD RN NET52 VDD P18 W=1.2U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.68U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.68U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=0.87U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NETQ VDD P18 W=1.2U L=0.18U
MN6 NETQ NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=1.12U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.12U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=1.1U PW=1.1U
XI21 NET80 SN IVG PW=0.81U NW=0.54U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSRHD1X                                                            *
* LAST TIME SAVED: MAR  4 16:19:08 2003                                       *
*******************************************************************************
.SUBCKT LATSRHD1X Q QN D G RN SN
MP8 VDD RN NET52 VDD P18 W=0.84U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.6U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.6U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NETQ VDD P18 W=0.84U L=0.18U
MN6 NETQ NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=1.06U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.06U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET80 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSHDLX                                                             *
* LAST TIME SAVED: MAR  4 16:18:52 2003                                       *
*******************************************************************************
.SUBCKT LATSHDLX Q QN D G SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.54U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.54U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1U L=0.18U
MN3 NET44 D GND GND N18 W=0.77U L=0.18U
MN6 NETQ NET73 GND GND N18 W=0.42U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSHD4X                                                             *
* LAST TIME SAVED: MAR  4 16:18:35 2003                                       *
*******************************************************************************
.SUBCKT LATSHD4X Q QN D G SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=3.36U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=3.36U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1.16U L=0.18U
MN3 NET44 D GND GND N18 W=1.86U L=0.18U
MN6 NETQ NET73 GND GND N18 W=0.6U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NETQ NET55 NET32 TG1G NW=1.18U PW=1.18U
XI21 NET73 SN IVG PW=1.05U NW=0.7U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSHD2X                                                             *
* LAST TIME SAVED: MAR  4 16:18:16 2003                                       *
*******************************************************************************
.SUBCKT LATSHD2X Q QN D G SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.68U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.68U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1.56U L=0.18U
MN3 NET44 D GND GND N18 W=0.9U L=0.18U
MN6 NETQ NET73 GND GND N18 W=0.72U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NETQ NET55 NET32 TG1G NW=1.1U PW=1.1U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATSHD1X                                                             *
* LAST TIME SAVED: MAR  4 16:18:00 2003                                       *
*******************************************************************************
.SUBCKT LATSHD1X Q QN D G SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.6U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.6U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1U L=0.18U
MN3 NET44 D GND GND N18 W=0.86U L=0.18U
MN6 NETQ NET73 GND GND N18 W=0.42U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATRHDLX                                                             *
* LAST TIME SAVED: MAR  4 16:17:40 2003                                       *
*******************************************************************************
.SUBCKT LATRHDLX Q QN D G RN
MP1 VDD D NET47 VDD P18 W=0.93U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NETQ VDD P18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=0.77U L=0.18U
MN2 NET47 D NET44 GND N18 W=0.77U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATRHD4X                                                             *
* LAST TIME SAVED: MAR  4 16:17:24 2003                                       *
*******************************************************************************
.SUBCKT LATRHD4X Q QN D G RN
MP1 VDD D NET47 VDD P18 W=3.44U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NETQ VDD P18 W=1.08U L=0.18U
MN3 NET44 RN GND GND N18 W=2.36U L=0.18U
MN2 NET47 D NET44 GND N18 W=2.36U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=1.18U PW=1.18U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATRHD2X                                                             *
* LAST TIME SAVED: MAR  4 16:17:08 2003                                       *
*******************************************************************************
.SUBCKT LATRHD2X Q QN D G RN
MP1 VDD D NET47 VDD P18 W=1.42U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NETQ VDD P18 W=1.08U L=0.18U
MN3 NET44 RN GND GND N18 W=1.18U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.18U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=1.1U PW=1.1U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATRHD1X                                                             *
* LAST TIME SAVED: MAR  4 16:16:52 2003                                       *
*******************************************************************************
.SUBCKT LATRHD1X Q QN D G RN
MP1 VDD D NET47 VDD P18 W=1.28U L=0.18U
MP4 NET26 NET55 NETQ VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NETQ VDD P18 W=0.6U L=0.18U
MN3 NET44 RN GND GND N18 W=1.06U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.06U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.3U L=0.18U
MN1 NETQ NET32 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NETQ NET55 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSRHDLX                                                           *
* LAST TIME SAVED: MAR  4 16:09:07 2003                                       *
*******************************************************************************
.SUBCKT LATNSRHDLX Q QN D GN RN SN
MP8 VDD RN NET52 VDD P18 W=0.84U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.16U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.16U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NET53 VDD P18 W=0.84U L=0.18U
MN6 NET53 NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=0.77U L=0.18U
MN2 NET47 D NET44 GND N18 W=0.77U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=0.7U PW=0.7U
XI21 NET80 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=0.64U NW=0.42U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSRHD4X                                                           *
* LAST TIME SAVED: MAR  4 16:08:52 2003                                       *
*******************************************************************************
.SUBCKT LATNSRHD4X Q QN D GN RN SN
MP8 VDD RN NET52 VDD P18 W=1.44U L=0.18U
MP6 NET103 D NET47 VDD P18 W=3.3U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=3.3U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1.68U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NET53 VDD P18 W=1.44U L=0.18U
MN6 NET53 NET80 GND GND N18 W=0.72U L=0.18U
MN3 NET44 RN GND GND N18 W=2.3U L=0.18U
MN2 NET47 D NET44 GND N18 W=2.3U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.8U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=1.18U PW=1.18U
XI21 NET80 SN IVG PW=1.5U NW=1U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NET53 IVG PW=4.8U NW=3.2U
XI10 NETQN NET53 IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSRHD2X                                                           *
* LAST TIME SAVED: MAR  4 16:08:34 2003                                       *
*******************************************************************************
.SUBCKT LATNSRHD2X Q QN D GN RN SN
MP8 VDD RN NET52 VDD P18 W=1.2U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.68U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.68U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=0.86U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NET53 VDD P18 W=1.2U L=0.18U
MN6 NET53 NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=1.12U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.12U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=1.1U PW=1.1U
XI21 NET80 SN IVG PW=0.81U NW=0.54U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NET53 IVG PW=2.4U NW=1.6U
XI10 NETQN NET53 IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSRHD1X                                                           *
* LAST TIME SAVED: MAR  4 16:08:17 2003                                       *
*******************************************************************************
.SUBCKT LATNSRHD1X Q QN D GN RN SN
MP8 VDD RN NET52 VDD P18 W=0.84U L=0.18U
MP6 NET103 D NET47 VDD P18 W=1.6U L=0.18U
MP1 VDD NET80 NET103 VDD P18 W=1.6U L=0.18U
MP7 VDD NET80 NET112 VDD P18 W=1U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.45U L=0.18U
MP5 NET112 NETQN NET26 VDD P18 W=0.45U L=0.18U
MP3 NET52 NET80 NET53 VDD P18 W=0.84U L=0.18U
MN6 NET53 NET80 GND GND N18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=1.06U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.06U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=0.7U PW=0.7U
XI21 NET80 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=1.2U NW=0.8U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSHDLX                                                            *
* LAST TIME SAVED: MAR  4 16:04:00 2003                                       *
*******************************************************************************
.SUBCKT LATNSHDLX Q QN D GN SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.54U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.54U L=0.18U
MP4 NET26 NET82 NET53 VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1U L=0.18U
MN3 NET44 D GND GND N18 W=0.77U L=0.18U
MN6 NET53 NET73 GND GND N18 W=0.42U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET32 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NET53 NET82 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET32 NET82 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=0.64U NW=0.42U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET82 GN IVG PW=0.84U NW=0.42U
.ENDS LATNSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSHD4X                                                            *
* LAST TIME SAVED: MAR 13 12:42:45 2003                                       *
*******************************************************************************
.SUBCKT LATNSHD4X Q QN D GN SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=3.36U L=0.18U
MP1 VDD NET61 NET47 VDD P18 W=3.36U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.6U L=0.18U
MP5 VDD NET61 NET48 VDD P18 W=1.64U L=0.18U
MN3 NET44 D GND GND N18 W=1.86U L=0.18U
MN6 NET53 NET61 GND GND N18 W=0.72U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET55 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NET53 NET32 NET55 TG1G NW=1.18U PW=1.18U
XI21 NET61 SN IVG PW=1.05U NW=0.7U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NET53 IVG PW=4.8U NW=3.2U
XI10 NETQN NET53 IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSHD2X                                                            *
* LAST TIME SAVED: MAR  4 16:03:31 2003                                       *
*******************************************************************************
.SUBCKT LATNSHD2X Q QN D GN SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.68U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.68U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1.68U L=0.18U
MN3 NET44 D GND GND N18 W=0.9U L=0.18U
MN6 NET53 NET73 GND GND N18 W=0.72U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET55 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NET53 NET32 NET55 TG1G NW=1.1U PW=1.1U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NET53 IVG PW=2.4U NW=1.6U
XI10 NETQN NET53 IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNSHD1X                                                            *
* LAST TIME SAVED: MAR  4 16:03:12 2003                                       *
*******************************************************************************
.SUBCKT LATNSHD1X Q QN D GN SN
MP7 NET48 NETQN NET26 VDD P18 W=0.6U L=0.18U
MP6 NET47 D NET44 VDD P18 W=1.6U L=0.18U
MP1 VDD NET73 NET47 VDD P18 W=1.6U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.6U L=0.18U
MP5 VDD NET73 NET48 VDD P18 W=1U L=0.18U
MN3 NET44 D GND GND N18 W=0.86U L=0.18U
MN6 NET53 NET73 GND GND N18 W=0.42U L=0.18U
MN5 NET38 NETQN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET55 NET38 GND N18 W=0.3U L=0.18U
XI9 NET44 NET53 NET32 NET55 TG1G NW=0.7U PW=0.7U
XI21 NET73 SN IVG PW=0.64U NW=0.42U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=1.2U NW=0.8U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNRHDLX                                                            *
* LAST TIME SAVED: MAR  4 16:02:55 2003                                       *
*******************************************************************************
.SUBCKT LATNRHDLX Q QN D GN RN
MP1 VDD D NET47 VDD P18 W=0.93U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NET53 VDD P18 W=0.42U L=0.18U
MN3 NET44 RN GND GND N18 W=0.77U L=0.18U
MN2 NET47 D NET44 GND N18 W=0.77U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET72 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET72 TG1G NW=0.7U PW=0.7U
XI13 NET72 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=0.64U NW=0.42U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNRHD4X                                                            *
* LAST TIME SAVED: MAR  4 16:02:38 2003                                       *
*******************************************************************************
.SUBCKT LATNRHD4X Q QN D GN RN
MP1 VDD D NET47 VDD P18 W=3.44U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NET53 VDD P18 W=1.08U L=0.18U
MN3 NET44 RN GND GND N18 W=2.36U L=0.18U
MN2 NET47 D NET44 GND N18 W=2.36U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=1.18U PW=1.18U
XI13 NET55 NET32 IVG PW=0.96U NW=0.48U
XI12 Q NET53 IVG PW=4.8U NW=3.2U
XI10 NETQN NET53 IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNRHD2X                                                            *
* LAST TIME SAVED: MAR  4 16:02:19 2003                                       *
*******************************************************************************
.SUBCKT LATNRHD2X Q QN D GN RN
MP1 VDD D NET47 VDD P18 W=1.42U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NET53 VDD P18 W=1.08U L=0.18U
MN3 NET44 RN GND GND N18 W=1.12U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.12U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=1.1U PW=1.1U
XI13 NET55 NET32 IVG PW=0.84U NW=0.42U
XI12 Q NET53 IVG PW=2.4U NW=1.6U
XI10 NETQN NET53 IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNRHD1X                                                            *
* LAST TIME SAVED: MAR  4 16:02:04 2003                                       *
*******************************************************************************
.SUBCKT LATNRHD1X Q QN D GN RN
MP1 VDD D NET47 VDD P18 W=1.28U L=0.18U
MP4 NET26 NET32 NET53 VDD P18 W=0.36U L=0.18U
MP5 VDD NETQN NET26 VDD P18 W=0.36U L=0.18U
MP3 VDD RN NET53 VDD P18 W=0.6U L=0.18U
MN3 NET44 RN GND GND N18 W=1.06U L=0.18U
MN2 NET47 D NET44 GND N18 W=1.06U L=0.18U
MN4 NET41 NETQN NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 RN GND GND N18 W=0.3U L=0.18U
MN1 NET53 NET55 NET41 GND N18 W=0.3U L=0.18U
XI9 NET47 NET53 NET32 NET55 TG1G NW=0.7U PW=0.7U
XI13 NET55 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET53 IVG PW=1.2U NW=0.8U
XI10 NETQN NET53 IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNHDLX                                                             *
* LAST TIME SAVED: MAR  4 16:01:45 2003                                       *
*******************************************************************************
.SUBCKT LATNHDLX Q QN D GN
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET32 NET24 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNHD4X                                                             *
* LAST TIME SAVED: MAR  4 16:01:31 2003                                       *
*******************************************************************************
.SUBCKT LATNHD4X Q QN D GN
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET32 NET24 TG1G NW=1.18U PW=1.18U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNHD2X                                                             *
* LAST TIME SAVED: MAR  4 16:01:14 2003                                       *
*******************************************************************************
.SUBCKT LATNHD2X Q QN D GN
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET32 NET24 TG1G NW=1.1U PW=1.1U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 GN IVG PW=1.2U NW=0.6U
.ENDS LATNHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATNHD1X                                                             *
* LAST TIME SAVED: MAR  4 16:00:50 2003                                       *
*******************************************************************************
.SUBCKT LATNHD1X Q QN D GN
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQ NET32 NET24 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 GN IVG PW=0.84U NW=0.42U
.ENDS LATNHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATHDLX                                                              *
* LAST TIME SAVED: MAR  4 16:00:33 2003                                       *
*******************************************************************************
.SUBCKT LATHDLX Q QN D G
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=0.64U NW=0.42U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATHD4X                                                              *
* LAST TIME SAVED: MAR  4 16:00:17 2003                                       *
*******************************************************************************
.SUBCKT LATHD4X Q QN D G
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQN NET24 NET32 TG1G NW=1.18U PW=1.18U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI12 QN NETQN IVG PW=4.8U NW=3.2U
XI10 NETQ NETQN IVG PW=1.68U NW=1.14U
XI5 Q NETQ IVG PW=4.8U NW=3.2U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATHD2XSPG                                                           *
* LAST TIME SAVED: MAR  4 16:00:00 2003                                       *
*******************************************************************************
.SUBCKT LATHD2XSPG Q QN D G
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATHD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATHD2X                                                              *
* LAST TIME SAVED: MAR  4 15:59:43 2003                                       *
*******************************************************************************
.SUBCKT LATHD2X Q QN D G
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 G IVG PW=1.2U NW=0.6U
.ENDS LATHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LATHD1X                                                              *
* LAST TIME SAVED: MAR  4 15:59:27 2003                                       *
*******************************************************************************
.SUBCKT LATHD1X Q QN D G
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 D NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=1.2U NW=0.8U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET32 G IVG PW=0.84U NW=0.42U
.ENDS LATHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHDLX                                                            *
* LAST TIME SAVED: AUG 30 10:45:03 2002                                       *
*******************************************************************************
.SUBCKT INVTSHDLX Z A E
MP0 VDD A NET9 VDD P18 W=1.2U L=0.18U
MP1 NET9 NET17 Z VDD P18 W=1.2U L=0.18U
MN1 NET12 A GND GND N18 W=0.8U L=0.18U
MN0 Z E NET12 GND N18 W=0.8U L=0.18U
XI0 NET17 E IVG PW=0.42U NW=0.3U
.ENDS INVTSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD8X                                                            *
* LAST TIME SAVED: AUG 30 10:44:58 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD8X Z A E
MN0 Z NET9 GND GND N18 W=6.4U L=0.18U
MN1 NET9 NET27 GND GND N18 W=2.4U L=0.18U
MN2 NET9 NET29 GND GND N18 W=0.8U L=0.18U
MP0 VDD NET27 NET14 VDD P18 W=3.44U L=0.18U
MP1 VDD E NET14 VDD P18 W=1.2U L=0.18U
MP4 VDD NET14 Z VDD P18 W=9.6U L=0.18U
XI6 NET9 NET14 E NET29 TG1G NW=1.2U PW=1.72U
XI7 NET27 A IVG PW=1.14U NW=0.76U
XI3 NET29 E IVG PW=0.48U NW=0.32U
.ENDS INVTSHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD4X                                                            *
* LAST TIME SAVED: AUG 30 10:44:53 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD4X Z A E
XI3 NET5 E IVG PW=0.42U NW=0.30U
XI7 NET7 A IVG PW=0.56U NW=0.38U
XI6 NET26 NET19 E NET5 TG1G NW=0.7U PW=0.7U
MP4 VDD NET19 Z VDD P18 W=4.8U L=0.18U
MP1 VDD E NET19 VDD P18 W=0.6U L=0.18U
MP0 VDD NET7 NET19 VDD P18 W=1.72U L=0.18U
MN2 NET26 NET5 GND GND N18 W=0.42U L=0.18U
MN1 NET26 NET7 GND GND N18 W=1.2U L=0.18U
MN0 Z NET26 GND GND N18 W=3.2U L=0.18U
.ENDS INVTSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD3X                                                            *
* LAST TIME SAVED: AUG 30 10:44:50 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD3X Z A E
MN2 NET9 NET29 GND GND N18 W=0.42U L=0.18U
MN1 NET9 NET27 GND GND N18 W=0.96U L=0.18U
MN0 Z NET9 GND GND N18 W=2.4U L=0.18U
MP4 VDD NET14 Z VDD P18 W=3.6U L=0.18U
MP1 VDD E NET14 VDD P18 W=0.64U L=0.18U
MP0 VDD NET27 NET14 VDD P18 W=1.44U L=0.18U
XI6 NET9 NET14 E NET29 TG1G NW=0.6U PW=0.6U
XI3 NET29 E IVG PW=0.45U NW=0.30U
XI7 NET27 A IVG PW=0.45U NW=0.30U
.ENDS INVTSHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD2X                                                            *
* LAST TIME SAVED: AUG 30 10:44:46 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD2X Z A E
MP0 VDD A NET9 VDD P18 W=4.8U L=0.18U
MP1 NET9 NET17 Z VDD P18 W=4.8U L=0.18U
MN0 Z E NET15 GND N18 W=3.2U L=0.18U
MN1 NET15 A GND GND N18 W=3.2U L=0.18U
XI0 NET17 E IVG PW=0.9U NW=0.6U
.ENDS INVTSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD20X                                                           *
* LAST TIME SAVED: AUG 30 10:44:49 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD20X Z A E
XI3 NET5 E IVG PW=1.2U NW=0.8U
XI7 NET7 A IVG PW=2.88U NW=1.82U
XI6 NET26 NET19 E NET5 TG1G NW=3.5U PW=3.5U
MP4 VDD NET19 Z VDD P18 W=24U L=0.18U
MP1 VDD E NET19 VDD P18 W=2.84U L=0.18U
MP0 VDD NET7 NET19 VDD P18 W=8.4U L=0.18U
MN2 NET26 NET5 GND GND N18 W=2.0U L=0.18U
MN1 NET26 NET7 GND GND N18 W=5.6U L=0.18U
MN0 Z NET26 GND GND N18 W=16U L=0.18U
.ENDS INVTSHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD1X                                                            *
* LAST TIME SAVED: AUG 30 10:44:41 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD1X Z A E
XI0 NET32 E IVG PW=0.45U NW=0.3U
MN0 Z E NET6 GND N18 W=1.6U L=0.18U
MN1 NET6 A GND GND N18 W=1.6U L=0.18U
MP1 NET12 NET32 Z VDD P18 W=2.4U L=0.18U
MP0 VDD A NET12 VDD P18 W=2.4U L=0.18U
.ENDS INVTSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD16X                                                           *
* LAST TIME SAVED: AUG 30 10:44:45 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD16X Z A E
MN0 Z NET9 GND GND N18 W=12.8U L=0.18U
MN1 NET9 NET27 GND GND N18 W=4.8U L=0.18U
MN2 NET9 NET29 GND GND N18 W=1.6U L=0.18U
MP0 VDD NET27 NET14 VDD P18 W=6.88U L=0.18U
MP1 VDD E NET14 VDD P18 W=2.4U L=0.18U
MP4 VDD NET14 Z VDD P18 W=19.2U L=0.18U
XI6 NET9 NET14 E NET29 TG1G NW=2.36U PW=2.36U
XI7 NET27 A IVG PW=2.24U NW=1.5U
XI3 NET29 E IVG PW=0.96U NW=0.64U
.ENDS INVTSHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVTSHD12X                                                           *
* LAST TIME SAVED: AUG 30 10:44:42 2002                                       *
*******************************************************************************
.SUBCKT INVTSHD12X Z A E
XI3 NET5 E IVG PW=0.72U NW=0.48U
XI7 NET7 A IVG PW=1.72U NW=1.14U
XI6 NET26 NET19 E NET5 TG1G NW=1.8U PW=1.8U
MP4 VDD NET19 Z VDD P18 W=14.4U L=0.18U
MP1 VDD E NET19 VDD P18 W=1.72U L=0.18U
MP0 VDD NET7 NET19 VDD P18 W=4.8U L=0.18U
MN2 NET26 NET5 GND GND N18 W=1.2U L=0.18U
MN1 NET26 NET7 GND GND N18 W=3.2U L=0.18U
MN0 Z NET26 GND GND N18 W=9.6U L=0.18U
.ENDS INVTSHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVODHD8X                                                            *
* LAST TIME SAVED: DEC 27 23:00:59 2003                                       *
*******************************************************************************
.SUBCKT INVODHD8X Z0 Z1 Z2 Z3 Z4 Z5 Z6 Z7 A
MN14 Z7 NET35 GND GND N18 W=1.6U L=0.18U
MN13 Z6 NET35 GND GND N18 W=1.6U L=0.18U
MN12 Z5 NET35 GND GND N18 W=1.6U L=0.18U
MN11 Z4 NET35 GND GND N18 W=1.6U L=0.18U
MN10 Z3 NET35 GND GND N18 W=1.6U L=0.18U
MN9 Z2 NET35 GND GND N18 W=1.6U L=0.19U
MN8 Z1 NET35 GND GND N18 W=1.6U L=0.19U
MN0 Z0 NET35 GND GND N18 W=1.6U L=0.18U
XI0 NET35 A IVG PW=2.4U NW=1.6U
.ENDS INVODHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHDPX                                                              *
* LAST TIME SAVED: AUG 30 10:34:57 2002                                       *
*******************************************************************************
.SUBCKT INVHDPX Z A
XI0 Z A IVG PW=1.72U NW=1.2U
.ENDS INVHDPX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHDLX                                                              *
* LAST TIME SAVED: AUG 30 10:34:55 2002                                       *
*******************************************************************************
.SUBCKT INVHDLX Z A
XI0 Z A IVG PW=0.64U NW=0.42U
.ENDS INVHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD8X                                                              *
* LAST TIME SAVED: AUG 30 10:34:52 2002                                       *
*******************************************************************************
.SUBCKT INVHD8X Z A
XI0 Z A IVG PW=9.6U NW=6.4U
.ENDS INVHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD4X                                                              *
* LAST TIME SAVED: AUG 30 10:34:50 2002                                       *
*******************************************************************************
.SUBCKT INVHD4X Z A
XI0 Z A IVG PW=4.8U NW=3.2U
.ENDS INVHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD3X                                                              *
* LAST TIME SAVED: AUG 30 10:34:48 2002                                       *
*******************************************************************************
.SUBCKT INVHD3X Z A
XI0 Z A IVG PW=3.6U NW=2.4U
.ENDS INVHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD2XSPG                                                           *
* LAST TIME SAVED: AUG 30 10:34:47 2002                                       *
*******************************************************************************
.SUBCKT INVHD2XSPG Z A
XI0 Z A IVG PW=2.4U NW=1.6U
.ENDS INVHD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD2X                                                              *
* LAST TIME SAVED: AUG 30 10:34:44 2002                                       *
*******************************************************************************
.SUBCKT INVHD2X Z A
XI0 Z A IVG PW=2.4U NW=1.6U
.ENDS INVHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD20X                                                             *
* LAST TIME SAVED: AUG 30 10:34:46 2002                                       *
*******************************************************************************
.SUBCKT INVHD20X Z A
XI0 Z NET8 IVG PW=24U NW=16U
XI1 NET6 A IVG PW=2U NW=1.2U
XI2 NET8 NET6 IVG PW=6U NW=4U
.ENDS INVHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD1X                                                              *
* LAST TIME SAVED: AUG 30 10:34:38 2002                                       *
*******************************************************************************
.SUBCKT INVHD1X Z A
XI0 Z A IVG PW=1.2U NW=0.77U
.ENDS INVHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD16X                                                             *
* LAST TIME SAVED: AUG 30 10:34:42 2002                                       *
*******************************************************************************
.SUBCKT INVHD16X Z A
XI0 Z NET8 IVG PW=19.2U NW=12.8U
XI1 NET6 A IVG PW=1.6U NW=1.1U
XI2 NET8 NET6 IVG PW=4.8U NW=3.2U
.ENDS INVHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVHD12X                                                             *
* LAST TIME SAVED: AUG 30 10:34:40 2002                                       *
*******************************************************************************
.SUBCKT INVHD12X Z A
XI2 NET4 NET6 IVG PW=3.6U NW=2.4U
XI1 NET6 A IVG PW=1.2U NW=0.8U
XI0 Z NET4 IVG PW=14.4U NW=9.6U
.ENDS INVHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHDLX                                                           *
* LAST TIME SAVED: AUG 30 10:32:34 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHDLX Z A
XI0 Z A IVG PW=0.96U NW=0.3U
.ENDS INVCLKHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD8X                                                           *
* LAST TIME SAVED: AUG 30 10:32:31 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD8X Z A
XI0 Z A IVG PW=9.6U NW=4.0U
.ENDS INVCLKHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD80X                                                          *
* LAST TIME SAVED: AUG 30 10:32:32 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD80X Z A
XI1 NET8 A IVG PW=6U NW=4.4U
XI2 NET6 NET8 IVG PW=24U NW=12U
XI0 Z NET6 IVG PW=96U NW=40U
.ENDS INVCLKHD80X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD4X                                                           *
* LAST TIME SAVED: AUG 30 10:32:27 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD4X Z A
XI0 Z A IVG PW=4.8U NW=1.92U
.ENDS INVCLKHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD40X                                                          *
* LAST TIME SAVED: AUG 30 10:32:29 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD40X Z A
XI1 NET8 A IVG PW=3U NW=2.2U
XI2 NET6 NET8 IVG PW=12U NW=6U
XI0 Z NET6 IVG PW=48U NW=19U
.ENDS INVCLKHD40X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD3X                                                           *
* LAST TIME SAVED: AUG 30 10:32:23 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD3X Z A
XI0 Z A IVG PW=3.6U NW=1.44U
.ENDS INVCLKHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD30X                                                          *
* LAST TIME SAVED: AUG 30 10:32:25 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD30X Z A
XI1 NET8 A IVG PW=2U NW=1.2U
XI2 NET6 NET8 IVG PW=8U NW=5.8U
XI0 Z NET6 IVG PW=36U NW=16.4U
.ENDS INVCLKHD30X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD2X                                                           *
* LAST TIME SAVED: AUG 30 10:32:20 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD2X Z A
XI0 Z A IVG PW=2.4U NW=0.94U
.ENDS INVCLKHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD20X                                                          *
* LAST TIME SAVED: AUG 30 10:32:21 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD20X Z A
XI0 Z A IVG PW=24U NW=10.3U
.ENDS INVCLKHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD1X                                                           *
* LAST TIME SAVED: AUG 30 10:32:10 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD1X Z A
XI0 Z A IVG PW=1.2U NW=0.4U
.ENDS INVCLKHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD16X                                                          *
* LAST TIME SAVED: AUG 30 10:32:18 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD16X Z A
XI0 Z A IVG PW=19.2U NW=8.2U
.ENDS INVCLKHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: INVCLKHD12X                                                          *
* LAST TIME SAVED: AUG 30 10:32:14 2002                                       *
*******************************************************************************
.SUBCKT INVCLKHD12X Z A
XI0 Z A IVG PW=14.4U NW=6.2U
.ENDS INVCLKHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: HOLDHD                                                               *
* LAST TIME SAVED: AUG 30 10:34:34 2002                                       *
*******************************************************************************
.SUBCKT HOLDHD Z
MN3 Z NET22 NET17 GND N18 W=0.3U L=0.36U
MN2 NET17 NET22 GND GND N18 W=0.3U L=0.36U
MP1 VDD NET22 Z VDD P18 W=0.3U L=0.36U
XI4 NET22 Z IVG PW=0.45U NW=0.3U
.ENDS HOLDHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: HAHDLX                                                               *
* LAST TIME SAVED: AUG 30 10:29:49 2002                                       *
*******************************************************************************
.SUBCKT HAHDLX CO S A B
XI1 NET_7 B A ND2G PW=0.51U NW=0.42U
XI3 NET45 NET_25 NET_23 B TG1G NW=0.6U PW=0.6U
XI4 A NET_25 B NET_23 TG1G NW=0.6U PW=0.6U
XI6 S NET_25 IVG PW=0.64U NW=0.42U
XI5 NET45 A IVG PW=0.64U NW=0.42U
XI2 CO NET_7 IVG PW=0.64U NW=0.42U
XI0 NET_23 B IVG PW=0.45U NW=0.3U
.ENDS HAHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: HAHD4X                                                               *
* LAST TIME SAVED: AUG 30 10:29:48 2002                                       *
*******************************************************************************
.SUBCKT HAHD4X CO S A B
XI1 NET_7 B A ND2G PW=1.72U NW=1.1U
XI3 NET45 NET_25 NET_21 B TG1G NW=2.0U PW=2.0U
XI4 A NET_25 B NET_21 TG1G NW=1.8U PW=1.8U
XI6 S NET_25 IVG PW=4.8U NW=3.2U
XI5 NET45 A IVG PW=3.6U NW=2.4U
XI2 CO NET_7 IVG PW=4.8U NW=3.2U
XI0 NET_21 B IVG PW=2.88U NW=1.92U
.ENDS HAHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: HAHD2X                                                               *
* LAST TIME SAVED: DEC 27 23:32:00 2003                                       *
*******************************************************************************
.SUBCKT HAHD2X CO S A B
XI7 S NET_57 IVG PW=2.4U NW=1.6U
XI0 NET_8 B IVG PW=1.44U NL=0.19U NW=0.96U
XI2 CO NET_23 IVG PW=2.4U NW=1.6U
XI5 NET45 A IVG PW=2.4U NW=1.6U
XI4 A NET_57 B NET_8 TG1G NW=1.0U PW=1.0U
XI3 NET45 NET_57 NET_8 B TG1G NW=1.2U PW=1.2U
XI1 NET_23 B A ND2G PW=1U NW=0.84U
.ENDS HAHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: HAHD1X                                                               *
* LAST TIME SAVED: AUG 30 10:29:44 2002                                       *
*******************************************************************************
.SUBCKT HAHD1X CO S A B
XI1 NET_7 B A ND2G PW=0.51U NW=0.42U
XI3 NET45 NET_25 NET_23 B TG1G NW=1U PW=1U
XI4 A NET_25 B NET_23 TG1G NW=0.8U PW=0.8U
XI6 S NET_25 IVG PW=1.2U NW=0.8U
XI5 NET45 A IVG PW=1.72U NW=1.2U
XI2 CO NET_7 IVG PW=1.2U NW=0.8U
XI0 NET_23 B IVG PW=0.72U NW=0.48U
.ENDS HAHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC8HD                                                           *
* LAST TIME SAVED: AUG 30 10:53:12 2002                                       *
*******************************************************************************
.SUBCKT FILLERC8HD
MP1 VDD GND VDD VDD P18 W=10.08U L=0.77U
.ENDS FILLERC8HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC6HD                                                           *
* LAST TIME SAVED: AUG 30 10:52:42 2002                                       *
*******************************************************************************
.SUBCKT FILLERC6HD
MP1 VDD GND VDD VDD P18 W=6.8U L=0.76U
.ENDS FILLERC6HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC64HD                                                          *
* LAST TIME SAVED: AUG 30 13:31:23 2002                                       *
*******************************************************************************
.SUBCKT FILLERC64HD
MP1 VDD GND VDD VDD P18 W=70.24U L=1.38U
.ENDS FILLERC64HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC4HD                                                           *
* LAST TIME SAVED: AUG 30 10:52:13 2002                                       *
*******************************************************************************
.SUBCKT FILLERC4HD
MP1 VDD GND VDD VDD P18 W=1.75U L=1.57U
.ENDS FILLERC4HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC3HD                                                           *
* LAST TIME SAVED: AUG 30 10:51:44 2002                                       *
*******************************************************************************
.SUBCKT FILLERC3HD
MP1 VDD GND VDD VDD P18 W=1.75U L=0.93U
.ENDS FILLERC3HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC32HD                                                          *
* LAST TIME SAVED: AUG 30 10:54:09 2002                                       *
*******************************************************************************
.SUBCKT FILLERC32HD
MP1 VDD GND VDD VDD P18 W=33.22U L=1.42U
.ENDS FILLERC32HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC2HD                                                           *
* LAST TIME SAVED: AUG 30 10:51:10 2002                                       *
*******************************************************************************
.SUBCKT FILLERC2HD
MP1 VDD GND VDD VDD P18 W=1.75U L=0.3U
.ENDS FILLERC2HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC1HD                                                           *
* LAST TIME SAVED: AUG 30 10:50:40 2002                                       *
*******************************************************************************
.SUBCKT FILLERC1HD
.ENDS FILLERC1HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FILLERC16HD                                                          *
* LAST TIME SAVED: AUG 30 10:53:39 2002                                       *
*******************************************************************************
.SUBCKT FILLERC16HD
MP1 VDD GND VDD VDD P18 W=16.99U L=1.27U
.ENDS FILLERC16HD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSRHDLX                                                          *
* LAST TIME SAVED: MAR 13 15:08:31 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSRHDLX Q QN CK J K RN SN TE TI
XI33 NET142 NET112 NET140 NET147 TRIIVG NW=0.3U PW=0.42U
MP4 NET40 NETQ NET39 VDD P18 W=1.2U L=0.18U
MP5 VDD NET62 NET39 VDD P18 W=0.72U L=0.18U
MP2 VDD NET155 NET97 VDD P18 W=1.16U L=0.18U
MP0 NET79 NET140 NETQ VDD P18 W=0.45U L=0.18U
MP3 VDD K NET40 VDD P18 W=1.2U L=0.18U
MP1 NET85 NET155 NETQ VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET85 VDD P18 W=0.84U L=0.18U
MP6 NET91 NET116 NET79 VDD P18 W=0.45U L=0.18U
MP7 VDD NET155 NET91 VDD P18 W=1U L=0.18U
MP9 NET97 NET142 NET112 VDD P18 W=1.16U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.6U L=0.18U
MN5 NET103 RN GND GND N18 W=0.6U L=0.18U
MN6 NETQ NET155 GND GND N18 W=0.42U L=0.18U
MN0 NET109 RN GND GND N18 W=0.77U L=0.18U
MN4 NET112 NET142 NET109 GND N18 W=0.77U L=0.18U
MN7 NETQ NET147 NET118 GND N18 W=0.3U L=0.18U
MN8 NET118 NET116 NET103 GND N18 W=0.3U L=0.18U
MN2 NET52 K GND GND N18 W=0.6U L=0.18U
MN1 NET39 NET62 NET52 GND N18 W=0.6U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
XI27 TI NET104 TE NET115 TG1G NW=0.42U PW=0.42U
XI9 NET112 NETQ NET140 NET147 TG1G NW=0.7U PW=0.7U
XI26 NET39 NET104 NET115 TE TG1G NW=0.8U PW=0.8U
XI6 NET104 NET142 NET147 NET140 TG1G NW=0.42U PW=0.42U
XI20 NET115 TE IVG PW=0.64U NW=0.42U
XI4 NET147 CK IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET116 NETQ IVG PW=0.64U NW=0.42U
XI5 QN NET116 IVG PW=0.64U NW=0.42U
XI21 NET155 SN IVG PW=0.64U NW=0.42U
XI13 NET140 NET147 IVG PW=0.6U NW=0.3U
.ENDS FFSJKSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSRHD4X                                                          *
* LAST TIME SAVED: MAR 13 15:05:52 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSRHD4X Q QN CK J K RN SN TE TI
XI33 NET131 NET107 NET129 NET130 TRIIVG NW=0.3U PW=0.42U
MP4 NET109 NETQ NET45 VDD P18 W=2.4U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET109 VDD P18 W=2.4U L=0.18U
MP2 VDD NET156 NET74 VDD P18 W=3.3U L=0.18U
MP7 VDD NET156 NET71 VDD P18 W=1.68U L=0.18U
MP9 NET83 NET156 NETQ VDD P18 W=1.44U L=0.18U
MP0 NET80 NET129 NETQ VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET83 VDD P18 W=1.44U L=0.18U
MP6 NET74 NET131 NET107 VDD P18 W=3.3U L=0.18U
MP1 NET71 NET108 NET80 VDD P18 W=0.45U L=0.18U
MN2 NET55 K GND GND N18 W=1.18U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=1.18U L=0.18U
MN3 NET55 NETQ GND GND N18 W=1.18U L=0.18U
MN7 NET182 RN GND GND N18 W=2.3U L=0.18U
MN6 NETQ NET156 GND GND N18 W=0.72U L=0.18U
MN8 NET110 NET108 NET101 GND N18 W=0.3U L=0.18U
MN0 NET107 NET131 NET182 GND N18 W=2.3U L=0.18U
MN4 NETQ NET130 NET110 GND N18 W=0.3U L=0.18U
MN5 NET101 RN GND GND N18 W=0.8U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
XI27 TI NET105 TE NET116 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET105 NET116 TE TG1G NW=0.8U PW=0.8U
XI6 NET105 NET131 NET130 NET129 TG1G NW=0.8U PW=0.8U
XI9 NET107 NETQ NET129 NET130 TG1G NW=1.18U PW=1.18U
XI20 NET116 TE IVG PW=0.64U NW=0.42U
XI4 NET130 CK IVG PW=1.2U NW=0.6U
XI21 NET156 SN IVG PW=1.5U NW=1U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NET108 NETQ IVG PW=1.68U NW=1.14U
XI5 QN NET108 IVG PW=4.8U NW=3.2U
XI13 NET129 NET130 IVG PW=0.96U NW=0.48U
.ENDS FFSJKSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSRHD2X                                                          *
* LAST TIME SAVED: MAR 13 15:03:32 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSRHD2X Q QN CK J K RN SN TE TI
XI33 NET131 NET185 NET148 NET146 TRIIVG NW=0.3U PW=0.42U
MP9 VDD NET156 NET88 VDD P18 W=1.68U L=0.18U
MP1 NET86 NET108 NET71 VDD P18 W=0.45U L=0.18U
MP2 NET83 NET156 NETQ VDD P18 W=1.2U L=0.18U
MP8 VDD RN NET83 VDD P18 W=1.2U L=0.18U
MP6 NET88 NET131 NET185 VDD P18 W=1.68U L=0.18U
MP7 VDD NET156 NET86 VDD P18 W=0.86U L=0.18U
MP0 NET71 NET148 NETQ VDD P18 W=0.45U L=0.18U
MP4 NET109 NETQ NET45 VDD P18 W=1.66U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET109 VDD P18 W=1.66U L=0.18U
MN4 NET185 NET131 NET101 GND N18 W=1.12U L=0.18U
MN6 NETQ NET156 GND GND N18 W=0.42U L=0.18U
MN5 NET110 NET108 NET107 GND N18 W=0.3U L=0.18U
MN7 NET107 RN GND GND N18 W=0.6U L=0.18U
MN8 NETQ NET146 NET110 GND N18 W=0.3U L=0.18U
MN0 NET101 RN GND GND N18 W=1.12U L=0.18U
MN3 NET55 NETQ GND GND N18 W=0.9U L=0.18U
MN2 NET55 K GND GND N18 W=0.9U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=0.9U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
XI9 NET185 NETQ NET148 NET146 TG1G NW=1.1U PW=1.1U
XI27 TI NET105 TE NET116 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET105 NET116 TE TG1G NW=0.8U PW=0.8U
XI6 NET105 NET131 NET146 NET148 TG1G NW=0.42U PW=0.42U
XI21 NET156 SN IVG PW=0.81U NW=0.54U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NET108 NETQ IVG PW=0.84U NW=0.56U
XI5 QN NET108 IVG PW=2.4U NW=1.6U
XI36 NET148 NET146 IVG PW=0.84U NW=0.42U
XI20 NET116 TE IVG PW=0.64U NW=0.42U
XI4 NET146 CK IVG PW=1.2U NW=0.6U
.ENDS FFSJKSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSRHD1X                                                          *
* LAST TIME SAVED: MAR 13 14:59:05 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSRHD1X Q QN CK J K RN SN TE TI
XI34 NET130 NET182 NET128 NET145 TRIIVG NW=0.3U PW=0.42U
MP4 NET107 NETQ NET45 VDD P18 W=1.6U L=0.18U
MP5 VDD NET58 NET45 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET107 VDD P18 W=1.6U L=0.18U
MP6 NET76 NET155 NETQ VDD P18 W=0.84U L=0.18U
MP1 VDD NET155 NET70 VDD P18 W=1.6U L=0.18U
MP8 VDD RN NET76 VDD P18 W=0.84U L=0.18U
MP9 NET70 NET130 NET182 VDD P18 W=1.6U L=0.18U
MP0 NET82 NET104 NET79 VDD P18 W=0.45U L=0.18U
MP7 VDD NET155 NET82 VDD P18 W=1U L=0.18U
MP2 NET79 NET128 NETQ VDD P18 W=0.45U L=0.18U
MN3 NET55 NETQ GND GND N18 W=0.8U L=0.18U
MN0 NETQ NET145 NET106 GND N18 W=0.3U L=0.18U
MN6 NETQ NET155 GND GND N18 W=0.42U L=0.18U
MN7 NET109 RN GND GND N18 W=1.06U L=0.18U
MN4 NET106 NET104 NET103 GND N18 W=0.3U L=0.18U
MN5 NET103 RN GND GND N18 W=0.6U L=0.18U
MN2 NET55 K GND GND N18 W=0.8U L=0.18U
MN1 NET45 NET58 NET55 GND N18 W=0.8U L=0.18U
MN8 NET182 NET130 NET109 GND N18 W=1.06U L=0.18U
XI18 NET58 NETQ J ND2G PW=0.51U NW=0.42U
XI27 TI NET100 TE NET115 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET100 NET115 TE TG1G NW=0.8U PW=0.8U
XI6 NET100 NET130 NET145 NET128 TG1G NW=0.42U PW=0.42U
XI9 NET182 NETQ NET128 NET145 TG1G NW=0.7U PW=0.7U
XI20 NET115 TE IVG PW=0.64U NW=0.42U
XI4 NET145 CK IVG PW=0.84U NW=0.42U
XI21 NET155 SN IVG PW=0.64U NW=0.42U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NET104 NETQ IVG PW=0.64U NW=0.42U
XI13 NET128 NET145 IVG PW=0.6U NW=0.3U
XI5 QN NET104 IVG PW=1.2U NW=0.8U
.ENDS FFSJKSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSHDLX                                                           *
* LAST TIME SAVED: MAR 13 14:57:08 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSHDLX Q QN CK J K SN TE TI
XI32 NET118 NET100 NET116 NET133 TRIIVG NW=0.3U PW=0.42U
MP4 NET44 NETQ NET43 VDD P18 W=1.2U L=0.18U
MP6 NET76 NET118 NET100 VDD P18 W=1.54U L=0.18U
MP5 VDD NET65 NET43 VDD P18 W=0.72U L=0.18U
MP7 NET73 NET101 NET82 VDD P18 W=0.6U L=0.18U
MP3 VDD K NET44 VDD P18 W=1.2U L=0.18U
MP2 VDD NET135 NET73 VDD P18 W=1U L=0.18U
MP0 NET82 NET116 NETQ VDD P18 W=0.6U L=0.18U
MP1 VDD NET135 NET76 VDD P18 W=1.54U L=0.18U
MN0 NETQ NET133 NET103 GND N18 W=0.3U L=0.18U
MN3 NET53 NETQ GND GND N18 W=0.6U L=0.18U
MN5 NET103 NET101 GND GND N18 W=0.3U L=0.18U
MN4 NET100 NET118 GND GND N18 W=0.77U L=0.18U
MN6 NETQ NET135 GND GND N18 W=0.42U L=0.18U
MN2 NET53 K GND GND N18 W=0.6U L=0.18U
MN1 NET43 NET65 NET53 GND N18 W=0.6U L=0.18U
XI18 NET65 NETQ J ND2G PW=0.51U NW=0.42U
XI30 TI NET99 TE NET110 TG1G NW=0.42U PW=0.42U
XI31 NET43 NET99 NET110 TE TG1G NW=0.8U PW=0.8U
XI9 NET100 NETQ NET116 NET133 TG1G NW=0.7U PW=0.7U
XI6 NET99 NET118 NET133 NET116 TG1G NW=0.42U PW=0.42U
XI4 NET133 CK IVG PW=0.84U NW=0.42U
XI20 NET110 TE IVG PW=0.64U NW=0.42U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI21 NET135 SN IVG PW=0.64U NW=0.42U
XI5 QN NET101 IVG PW=0.64U NW=0.42U
XI13 NET116 NET133 IVG PW=0.6U NW=0.3U
XI10 NET101 NETQ IVG PW=0.64U NW=0.42U
.ENDS FFSJKSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSHD4X                                                           *
* LAST TIME SAVED: DEC 27 18:42:40 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSHD4X Q QN CK J K SN TE TI
XI32 NET118 NET66 NET116 NET133 TRIIVG NW=0.3U PW=0.42U
MP4 NET44 NETQ NET75 VDD P18 W=2.4U L=0.18U
MP2 VDD NET137 NET82 VDD P18 W=1.64U L=0.18U
MP5 VDD NET65 NET75 VDD P18 W=1.42U L=0.18U
MP0 NET73 NET116 NETQ VDD P18 W=0.6U L=0.18U
MP3 VDD K NET44 VDD P18 W=2.4U L=0.18U
MP1 VDD NET137 NET79 VDD P18 W=3.36U L=0.18U
MP7 NET82 NET98 NET73 VDD P18 W=0.6U L=0.18U
MP6 NET79 NET118 NET66 VDD P18 W=3.36U L=0.18U
MN4 NET66 NET118 GND GND N18 W=1.86U L=0.19U
MN3 NET53 NETQ GND GND N18 W=1.18U L=0.18U
MN0 NETQ NET133 NET100 GND N18 W=0.3U L=0.18U
MN5 NET100 NET98 GND GND N18 W=0.3U L=0.18U
MN6 NETQ NET137 GND GND N18 W=0.72U L=0.18U
MN2 NET53 K GND GND N18 W=1.18U L=0.18U
MN1 NET75 NET65 NET53 GND N18 W=1.18U L=0.18U
XI18 NET65 NETQ J ND2G PW=0.51U NW=0.42U
XI6 NET99 NET118 NET133 NET116 TG1G NW=0.8U PW=0.8U
XI30 TI NET99 TE NET110 TG1G NW=0.42U PW=0.42U
XI31 NET75 NET99 NET110 TE TG1G NW=0.8U PW=0.8U
XI9 NET66 NETQ NET116 NET133 TG1G NW=1.18U PW=1.18U
XI4 NET133 CK IVG PW=1.2U NW=0.6U
XI20 NET110 TE IVG PW=0.64U NW=0.42U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI13 NET116 NET133 IVG PW=0.96U NW=0.48U
XI21 NET137 SN IVG PW=1.05U NW=0.7U
XI5 QN NET98 IVG PW=4.8U NW=3.2U
XI10 NET98 NETQ IVG PW=1.68U NW=1.14U
.ENDS FFSJKSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSHD2X                                                           *
* LAST TIME SAVED: MAR 13 14:54:21 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSHD2X Q QN CK J K SN TE TI
XI32 NET116 NET95 NET114 NET131 TRIIVG NW=0.3U PW=0.42U
MP4 NET36 NETQ NET35 VDD P18 W=1.66U L=0.18U
MP5 VDD NET66 NET35 VDD P18 W=1.08U L=0.18U
MP6 NET71 NET116 NET95 VDD P18 W=1.68U L=0.18U
MP3 VDD K NET36 VDD P18 W=1.66U L=0.18U
MP2 VDD NET139 NET74 VDD P18 W=1.68U L=0.18U
MP1 VDD NET139 NET71 VDD P18 W=1.68U L=0.18U
MP0 NET77 NET114 NETQ VDD P18 W=0.6U L=0.18U
MP7 NET74 NET90 NET77 VDD P18 W=0.6U L=0.18U
MN3 NET48 NETQ GND GND N18 W=0.9U L=0.18U
MN0 NETQ NET131 NET92 GND N18 W=0.3U L=0.18U
MN6 NETQ NET139 GND GND N18 W=0.72U L=0.18U
MN4 NET95 NET116 GND GND N18 W=0.9U L=0.18U
MN5 NET92 NET90 GND GND N18 W=0.3U L=0.18U
MN2 NET48 K GND GND N18 W=0.9U L=0.18U
MN1 NET35 NET66 NET48 GND N18 W=0.9U L=0.18U
XI18 NET66 NETQ J ND2G PW=0.51U NW=0.42U
XI30 TI NET155 TE NET166 TG1G NW=0.42U PW=0.42U
XI31 NET35 NET155 NET166 TE TG1G NW=0.8U PW=0.8U
XI9 NET95 NETQ NET114 NET131 TG1G NW=1.1U PW=1.1U
XI6 NET155 NET116 NET131 NET114 TG1G NW=0.42U PW=0.42U
XI4 NET131 CK IVG PW=1.2U NW=0.6U
XI20 NET166 TE IVG PW=0.64U NW=0.42U
XI5 QN NET90 IVG PW=2.4U NW=1.6U
XI10 NET90 NETQ IVG PW=0.84U NW=0.56U
XI13 NET114 NET131 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI21 NET139 SN IVG PW=0.64U NW=0.42U
.ENDS FFSJKSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKSHD1X                                                           *
* LAST TIME SAVED: MAR 13 14:52:36 2003                                       *
*******************************************************************************
.SUBCKT FFSJKSHD1X Q QN CK J K SN TE TI
XI32 NET119 NET91 NET117 NET130 TRIIVG NW=0.3U PW=0.42U
MP4 NET43 NETQ NET42 VDD P18 W=1.6U L=0.18U
MP5 VDD NET64 NET42 VDD P18 W=0.96U L=0.18U
MP6 NET70 NET119 NET91 VDD P18 W=1.6U L=0.18U
MP3 VDD K NET43 VDD P18 W=1.6U L=0.18U
MP2 NET67 NET117 NETQ VDD P18 W=0.6U L=0.18U
MP1 VDD NET138 NET70 VDD P18 W=1.6U L=0.18U
MP0 VDD NET138 NET73 VDD P18 W=1U L=0.18U
MP7 NET73 NET92 NET67 VDD P18 W=0.6U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.8U L=0.18U
MN6 NETQ NET138 GND GND N18 W=0.42U L=0.18U
MN0 NETQ NET130 NET94 GND N18 W=0.3U L=0.18U
MN5 NET94 NET92 GND GND N18 W=0.3U L=0.18U
MN4 NET91 NET119 GND GND N18 W=0.86U L=0.18U
MN2 NET52 K GND GND N18 W=0.8U L=0.18U
MN1 NET42 NET64 NET52 GND N18 W=0.8U L=0.18U
XI18 NET64 NETQ J ND2G PW=0.51U NW=0.42U
XI30 TI NET96 TE NET107 TG1G NW=0.42U PW=0.42U
XI31 NET42 NET96 NET107 TE TG1G NW=0.8U PW=0.8U
XI6 NET96 NET119 NET130 NET117 TG1G NW=0.42U PW=0.42U
XI9 NET91 NETQ NET117 NET130 TG1G NW=0.7U PW=0.7U
XI4 NET130 CK IVG PW=0.84U NW=0.42U
XI20 NET107 TE IVG PW=0.64U NW=0.42U
XI13 NET117 NET130 IVG PW=0.6U NW=0.3U
XI10 NET92 NETQ IVG PW=0.64U NW=0.42U
XI5 QN NET92 IVG PW=1.2U NW=0.8U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI21 NET138 SN IVG PW=0.64U NW=0.42U
.ENDS FFSJKSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKRHDLX                                                           *
* LAST TIME SAVED: NOV 25 17:49:59 2003                                       *
*******************************************************************************
.SUBCKT FFSJKRHDLX Q QN CK J K RN TE TI
XI33 NET142 NET112 NET140 NET147 TRIIVG NW=0.3U PW=0.42U
MP4 NET40 NETQ NET39 VDD P18 W=1.2U L=0.18U
MP5 VDD NET62 NET39 VDD P18 W=0.72U L=0.18U
MP0 NET79 NET140 NETQ VDD P18 W=0.45U L=0.18U
MP3 VDD K NET40 VDD P18 W=1.2U L=0.18U
MP8 VDD RN NETQ VDD P18 W=0.64U L=0.18U
MP6 VDD NET116 NET79 VDD P18 W=0.45U L=0.18U
MP9 VDD NET142 NET112 VDD P18 W=0.88U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.6U L=0.18U
MN5 NET103 RN GND GND N18 W=0.6U L=0.18U
MN0 NET109 RN GND GND N18 W=0.77U L=0.18U
MN4 NET112 NET142 NET109 GND N18 W=0.77U L=0.18U
MN7 NETQ NET147 NET118 GND N18 W=0.3U L=0.18U
MN8 NET118 NET116 NET103 GND N18 W=0.3U L=0.18U
MN2 NET52 K GND GND N18 W=0.6U L=0.18U
MN1 NET39 NET62 NET52 GND N18 W=0.6U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
XI27 TI NET104 TE NET115 TG1G NW=0.42U PW=0.42U
XI9 NET112 NETQ NET140 NET147 TG1G NW=0.7U PW=0.7U
XI26 NET39 NET104 NET115 TE TG1G NW=0.8U PW=0.8U
XI6 NET104 NET142 NET147 NET140 TG1G NW=0.42U PW=0.42U
XI20 NET115 TE IVG PW=0.64U NW=0.42U
XI4 NET147 CK IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET116 NETQ IVG PW=0.42U NW=0.3U
XI5 QN NET116 IVG PW=0.64U NW=0.42U
XI13 NET140 NET147 IVG PW=0.6U NW=0.3U
.ENDS FFSJKRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKRHD4X                                                           *
* LAST TIME SAVED: NOV 25 17:48:03 2003                                       *
*******************************************************************************
.SUBCKT FFSJKRHD4X Q QN CK J K RN TE TI
XI33 NET131 NET107 NET129 NET130 TRIIVG NW=0.3U PW=0.42U
MP4 NET109 NET83 NET45 VDD P18 W=2.4U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET109 VDD P18 W=2.4U L=0.18U
MP0 NET80 NET129 NET83 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET83 VDD P18 W=1.1U L=0.18U
MP6 VDD NET131 NET107 VDD P18 W=2.52U L=0.18U
MP1 VDD NET108 NET80 VDD P18 W=0.45U L=0.18U
MN2 NET55 K GND GND N18 W=1.18U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=1.18U L=0.18U
MN3 NET55 NET83 GND GND N18 W=1.18U L=0.18U
MN7 NET182 RN GND GND N18 W=2.3U L=0.18U
MN8 NET110 NET108 NET101 GND N18 W=0.3U L=0.18U
MN0 NET107 NET131 NET182 GND N18 W=2.3U L=0.18U
MN4 NET83 NET130 NET110 GND N18 W=0.3U L=0.18U
MN5 NET101 RN GND GND N18 W=0.8U L=0.18U
XI18 NET62 NET83 J ND2G PW=0.51U NW=0.42U
XI27 TI NET105 TE NET116 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET105 NET116 TE TG1G NW=0.8U PW=0.8U
XI6 NET105 NET131 NET130 NET129 TG1G NW=0.8U PW=0.8U
XI9 NET107 NET83 NET129 NET130 TG1G NW=1.18U PW=1.18U
XI20 NET116 TE IVG PW=0.64U NW=0.42U
XI4 NET130 CK IVG PW=1.2U NW=0.6U
XI12 Q NET83 IVG PW=4.8U NW=3.2U
XI10 NET108 NET83 IVG PW=1.68U NW=1.14U
XI5 QN NET108 IVG PW=4.8U NW=3.2U
XI13 NET129 NET130 IVG PW=0.96U NW=0.48U
.ENDS FFSJKRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKRHD2X                                                           *
* LAST TIME SAVED: NOV 25 17:46:09 2003                                       *
*******************************************************************************
.SUBCKT FFSJKRHD2X Q QN CK J K RN TE TI
XI33 NET131 NET185 NET148 NET146 TRIIVG NW=0.3U PW=0.42U
MP1 VDD NET108 NET71 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET83 VDD P18 W=0.64U L=0.18U
MP6 VDD NET131 NET185 VDD P18 W=1.28U L=0.18U
MP0 NET71 NET148 NET83 VDD P18 W=0.45U L=0.18U
MP4 NET109 NET83 NET45 VDD P18 W=1.66U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET109 VDD P18 W=1.66U L=0.18U
MN4 NET185 NET131 NET101 GND N18 W=1.12U L=0.18U
MN5 NET110 NET108 NET107 GND N18 W=0.3U L=0.18U
MN7 NET107 RN GND GND N18 W=0.6U L=0.18U
MN8 NET83 NET146 NET110 GND N18 W=0.3U L=0.18U
MN0 NET101 RN GND GND N18 W=1.12U L=0.18U
MN3 NET55 NET83 GND GND N18 W=0.9U L=0.18U
MN2 NET55 K GND GND N18 W=0.9U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=0.9U L=0.18U
XI18 NET62 NET83 J ND2G PW=0.51U NW=0.42U
XI9 NET185 NET83 NET148 NET146 TG1G NW=1.1U PW=1.1U
XI27 TI NET105 TE NET116 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET105 NET116 TE TG1G NW=0.8U PW=0.8U
XI6 NET105 NET131 NET146 NET148 TG1G NW=0.42U PW=0.42U
XI12 Q NET83 IVG PW=2.4U NW=1.6U
XI10 NET108 NET83 IVG PW=0.84U NW=0.56U
XI5 QN NET108 IVG PW=2.4U NW=1.6U
XI36 NET148 NET146 IVG PW=0.84U NW=0.42U
XI20 NET116 TE IVG PW=0.64U NW=0.42U
XI4 NET146 CK IVG PW=1.2U NW=0.6U
.ENDS FFSJKRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKRHD1X                                                           *
* LAST TIME SAVED: NOV 13 16:59:16 2003                                       *
*******************************************************************************
.SUBCKT FFSJKRHD1X Q QN CK J K RN TE TI
XI34 NET130 NET182 NET128 NET145 TRIIVG NW=0.3U PW=0.42U
MP4 NET107 NET76 NET45 VDD P18 W=1.6U L=0.18U
MP5 VDD NET58 NET45 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET107 VDD P18 W=1.6U L=0.18U
MP8 VDD RN NET76 VDD P18 W=0.64U L=0.18U
MP9 VDD NET130 NET182 VDD P18 W=1.28U L=0.18U
MP0 VDD NET104 NET79 VDD P18 W=0.45U L=0.18U
MP2 NET79 NET128 NET76 VDD P18 W=0.45U L=0.18U
MN3 NET55 NET76 GND GND N18 W=0.8U L=0.18U
MN0 NET76 NET145 NET106 GND N18 W=0.3U L=0.18U
MN7 NET109 RN GND GND N18 W=1.06U L=0.18U
MN4 NET106 NET104 NET103 GND N18 W=0.3U L=0.18U
MN5 NET103 RN GND GND N18 W=0.6U L=0.18U
MN2 NET55 K GND GND N18 W=0.8U L=0.18U
MN1 NET45 NET58 NET55 GND N18 W=0.8U L=0.18U
MN8 NET182 NET130 NET109 GND N18 W=1.06U L=0.18U
XI18 NET58 NET76 J ND2G PW=0.51U NW=0.42U
XI27 TI NET100 TE NET115 TG1G NW=0.42U PW=0.42U
XI26 NET45 NET100 NET115 TE TG1G NW=0.8U PW=0.8U
XI6 NET100 NET130 NET145 NET128 TG1G NW=0.42U PW=0.42U
XI9 NET182 NET76 NET128 NET145 TG1G NW=0.7U PW=0.7U
XI20 NET115 TE IVG PW=0.64U NW=0.42U
XI4 NET145 CK IVG PW=0.84U NW=0.42U
XI12 Q NET76 IVG PW=1.2U NW=0.8U
XI10 NET104 NET76 IVG PW=0.64U NW=0.42U
XI13 NET128 NET145 IVG PW=0.6U NW=0.3U
XI5 QN NET104 IVG PW=1.2U NW=0.8U
.ENDS FFSJKRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKHDLX                                                            *
* LAST TIME SAVED: MAR  4 15:47:53 2003                                       *
*******************************************************************************
.SUBCKT FFSJKHDLX Q QN CK J K TE TI
MP4 NET34 NETQ NET100 VDD P18 W=1.2U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=0.72U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.2U L=0.18U
MN2 NET101 K GND GND N18 W=0.6U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.6U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.6U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.52U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI27 TI NET88 TE NET99 TG1G NW=0.42U PW=0.42U
XI26 NET100 NET88 NET99 TE TG1G NW=0.8U PW=0.8U
XI6 NET88 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=0.7U PW=0.7U
XI20 NET99 TE IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET32 NET96 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET96 CK IVG PW=0.84U NW=0.42U
.ENDS FFSJKHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKHD4X                                                            *
* LAST TIME SAVED: MAR  4 15:47:37 2003                                       *
*******************************************************************************
.SUBCKT FFSJKHD4X Q QN CK J K TE TI
MP4 NET34 NETQ NET100 VDD P18 W=2.4U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET34 VDD P18 W=2.4U L=0.18U
MN2 NET101 K GND GND N18 W=1.18U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=1.18U L=0.18U
MN3 NET101 NETQ GND GND N18 W=1.18U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI27 TI NET88 TE NET99 TG1G NW=0.42U PW=0.42U
XI26 NET100 NET88 NET99 TE TG1G NW=0.8U PW=0.8U
XI6 NET88 NET33 NET96 NET32 TG1G NW=0.8U PW=0.8U
XI9 NET46 NETQ NET32 NET96 TG1G NW=1.18U PW=1.18U
XI20 NET99 TE IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=3.44U NW=2.44U
XI13 NET32 NET96 IVG PW=0.96U NW=0.48U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET96 CK IVG PW=1.2U NW=0.6U
.ENDS FFSJKHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKHD2X                                                            *
* LAST TIME SAVED: MAR  4 15:47:18 2003                                       *
*******************************************************************************
.SUBCKT FFSJKHD2X Q QN CK J K TE TI
MP4 NET34 NETQ NET100 VDD P18 W=1.66U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.66U L=0.18U
MN2 NET101 K GND GND N18 W=0.9U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.9U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.9U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI27 TI NET88 TE NET99 TG1G NW=0.42U PW=0.42U
XI26 NET100 NET88 NET99 TE TG1G NW=0.8U PW=0.8U
XI6 NET88 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=1.1U PW=1.1U
XI20 NET99 TE IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI13 NET32 NET96 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET96 CK IVG PW=1.2U NW=0.6U
.ENDS FFSJKHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSJKHD1X                                                            *
* LAST TIME SAVED: MAR  4 15:47:01 2003                                       *
*******************************************************************************
.SUBCKT FFSJKHD1X Q QN CK J K TE TI
MP4 NET34 NETQ NET100 VDD P18 W=1.6U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.6U L=0.18U
MN2 NET101 K GND GND N18 W=0.8U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.8U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.8U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI27 TI NET89 TE NET116 TG1G NW=0.42U PW=0.42U
XI26 NET100 NET89 NET116 TE TG1G NW=0.8U PW=0.8U
XI6 NET89 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=0.7U PW=0.7U
XI20 NET116 TE IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET32 NET96 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET96 CK IVG PW=0.84U NW=0.42U
.ENDS FFSJKHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDQHDLX                                                           *
* LAST TIME SAVED: DEC  1 14:33:09 2003                                       *
*******************************************************************************
.SUBCKT FFSEDQHDLX Q CK D E TE TI
XI23 NET42 NETQN NET61 E TRIIVG NW=0.32U PW=0.48U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI24 NET42 D E NET61 TRIIVG NW=0.32U PW=0.48U
XI27 NET33 NET58 NET32 NET24 TRIIVG NW=0.32U PW=0.48U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.42U PW=0.42U
XI25 NET78 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI26 NET78 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSEDQHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDQHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:32:49 2003                                       *
*******************************************************************************
.SUBCKT FFSEDQHD4X Q CK D E TE TI
XI23 NET42 NETQN NET61 E TRIIVG NW=0.6U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI24 NET42 D E NET61 TRIIVG NW=0.6U PW=0.9U
XI27 NET33 NET58 NET32 NET24 TRIIVG NW=1U PW=1.17U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.6U PW=0.6U
XI25 NET78 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.81U NW=1.81U
XI26 NET78 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
.ENDS FFSEDQHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDQHD2X                                                           *
* LAST TIME SAVED: DEC  1 14:32:28 2003                                       *
*******************************************************************************
.SUBCKT FFSEDQHD2X Q CK D E TE TI
XI23 NET42 NETQN NET61 E TRIIVG NW=0.42U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI24 NET42 D E NET61 TRIIVG NW=0.42U PW=0.64U
XI27 NET33 NET58 NET32 NET24 TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.42U PW=0.42U
XI25 NET78 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI26 NET78 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFSEDQHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDQHD1X                                                           *
* LAST TIME SAVED: DEC  1 14:31:58 2003                                       *
*******************************************************************************
.SUBCKT FFSEDQHD1X Q CK D E TE TI
XI23 NET42 NETQN NET61 E TRIIVG NW=0.42U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI24 NET42 D E NET61 TRIIVG NW=0.42U PW=0.64U
XI27 NET33 NET58 NET32 NET24 TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.42U PW=0.42U
XI25 NET78 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI26 NET78 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSEDQHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDHDLX                                                            *
* LAST TIME SAVED: DEC  1 14:34:54 2003                                       *
*******************************************************************************
.SUBCKT FFSEDHDLX Q QN CK D E TE TI
XI24 NET42 D E NET61 TRIIVG NW=0.3U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET42 NETQ NET61 E TRIIVG NW=0.3U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.6U PW=0.6U
XI25 NET82 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.6U PW=0.6U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI26 NET82 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSEDHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:34:38 2003                                       *
*******************************************************************************
.SUBCKT FFSEDHD4X Q QN CK D E TE TI
XI24 NET42 D E NET61 TRIIVG NW=0.45U PW=1.62U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET42 NETQ NET61 E TRIIVG NW=0.45U PW=1.62U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=1.1U PW=1.1U
XI25 NET82 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=1.1U PW=1.1U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.52U NW=1.68U
XI26 NET82 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
.ENDS FFSEDHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDHD2X                                                            *
* LAST TIME SAVED: DEC  1 14:34:23 2003                                       *
*******************************************************************************
.SUBCKT FFSEDHD2X Q QN CK D E TE TI
XI24 NET42 D E NET61 TRIIVG NW=0.3U PW=1.05U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET42 NETQ NET61 E TRIIVG NW=0.3U PW=1.05U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.8U PW=0.8U
XI25 NET82 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.8U PW=0.8U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI26 NET82 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFSEDHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDHD1X                                                            *
* LAST TIME SAVED: DEC  1 14:34:06 2003                                       *
*******************************************************************************
.SUBCKT FFSEDHD1X Q QN CK D E TE TI
XI24 NET42 D E NET61 TRIIVG NW=0.3U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET42 NETQ NET61 E TRIIVG NW=0.3U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI21 NET42 NET58 NET81 TE TG1G NW=0.6U PW=0.6U
XI25 NET82 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.6U PW=0.6U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI22 NET81 TE IVG PW=0.42U NW=0.3U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI26 NET82 TI IVG PW=0.42U NW=0.3U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSEDHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDCRHDLX                                                          *
* LAST TIME SAVED: MAR  4 15:32:14 2003                                       *
*******************************************************************************
.SUBCKT FFSEDCRHDLX Q QN CK D E RN TE TI
XI18 NET63 RN NET54 ND2G PW=0.6U NW=0.5U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET63 NET58 NET81 TE TG1G NW=0.8U PW=0.8U
XI25 NET89 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI20 NETQN NET54 NET65 E TG1G NW=0.42U PW=0.42U
XI19 D NET54 E NET65 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI24 NET89 TI IVG PW=0.42U NW=0.3U
XI23 NET81 TE IVG PW=0.64U NW=0.42U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=0.64U NW=0.42U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFSEDCRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDCRHD4X                                                          *
* LAST TIME SAVED: MAR  4 15:31:55 2003                                       *
*******************************************************************************
.SUBCKT FFSEDCRHD4X Q QN CK D E RN TE TI
XI18 NET63 RN NET54 ND2G PW=1.47U NW=1.18U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI25 NET90 NET66 TE NET83 TG1G NW=0.42U PW=0.42U
XI22 NET63 NET66 NET83 TE TG1G NW=0.8U PW=0.8U
XI20 NETQN NET54 NET65 E TG1G NW=0.7U PW=0.7U
XI19 D NET54 E NET65 TG1G NW=0.7U PW=0.7U
XI6 NET66 NET33 NET32 NET24 TG1G NW=0.8U PW=0.8U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.18U PW=1.18U
XI24 NET90 TI IVG PW=0.42U NW=0.3U
XI23 NET83 TE IVG PW=0.64U NW=0.42U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=3.44U NW=2.3U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI12 QN NETQN IVG PW=4.8U NW=3.2U
XI10 NETQ NETQN IVG PW=1.68U NW=1.14U
XI5 Q NETQ IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFSEDCRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDCRHD2X                                                          *
* LAST TIME SAVED: MAR  4 15:31:37 2003                                       *
*******************************************************************************
.SUBCKT FFSEDCRHD2X Q QN CK D E RN TE TI
XI18 NET63 RN NET54 ND2G PW=0.96U NW=0.8U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET63 NET58 NET81 TE TG1G NW=0.8U PW=0.8U
XI20 NETQN NET54 NET65 E TG1G NW=0.6U PW=0.6U
XI19 D NET54 E NET65 TG1G NW=0.6U PW=0.6U
XI25 NET89 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI24 NET89 TI IVG PW=0.42U NW=0.3U
XI23 NET81 TE IVG PW=0.64U NW=0.42U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFSEDCRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSEDCRHD1X                                                          *
* LAST TIME SAVED: MAR  4 15:31:20 2003                                       *
*******************************************************************************
.SUBCKT FFSEDCRHD1X Q QN CK D E RN TE TI
XI18 NET63 RN NET54 ND2G PW=0.66U NW=0.55U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI25 NET91 NET58 TE NET81 TG1G NW=0.42U PW=0.42U
XI22 NET63 NET58 NET81 TE TG1G NW=0.8U PW=0.8U
XI20 NETQN NET54 NET65 E TG1G NW=0.6U PW=0.6U
XI19 D NET54 E NET65 TG1G NW=0.6U PW=0.6U
XI6 NET58 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI23 NET81 TE IVG PW=0.64U NW=0.42U
XI24 NET91 TI IVG PW=0.42U NW=0.3U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=1.2U NW=0.8U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFSEDCRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSRHDLX                                                           *
* LAST TIME SAVED: DEC  1 14:36:03 2003                                       *
*******************************************************************************
.SUBCKT FFSDSRHDLX Q QN CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.1U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.1U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.18U
MN0 NET55 SN NET180 GND N18 W=0.54U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET180 NET117 GND GND N18 W=0.54U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=0.72U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=0.72U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.5U PW=0.5U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=0.64U NW=0.32U
XI5 Q NET80 IVG PW=0.64U NW=0.32U
XI13 NET94 NET115 IVG PW=0.42U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSRHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:35:48 2003                                       *
*******************************************************************************
.SUBCKT FFSDSRHD4X Q QN CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=1.1U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=3.3U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=3.3U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1.68U L=0.18U
MN0 NET55 SN NET180 GND N18 W=0.92U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET180 NET117 GND GND N18 W=0.92U L=0.18U
MN5 NET142 SN GND GND N18 W=0.8U L=0.18U
MN3 NET73 SN GND GND N18 W=2.16U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=2.16U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG_1 NW=0.9U PW=1.5U PL0=0.19U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.7U PW=0.7U
XI21 NET117 RN IVG PW=1.5U NW=1.1U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.8U
XI12 QN NET55 IVG PW=4.8U NW=3.2U
XI5 Q NET80 IVG PW=4.8U NW=3.2U
XI13 NET94 NET115 IVG PW=0.93U NW=0.3U
XI10 NET80 NET55 IVG PW=1.77U NW=1.18U
.ENDS FFSDSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSRHD2X                                                           *
* LAST TIME SAVED: DEC  1 14:35:33 2003                                       *
*******************************************************************************
.SUBCKT FFSDSRHD2X Q QN CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=2.25U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=2.25U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=0.86U L=0.18U
MN0 NET55 SN NET180 GND N18 W=0.54U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET180 NET117 GND GND N18 W=0.54U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=1.57U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.57U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.1U PW=1.1U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.81U NW=0.54U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.45U
XI12 QN NET55 IVG PW=2.4U NW=1.6U
XI5 Q NET80 IVG PW=2.4U NW=1.6U
XI13 NET94 NET115 IVG PW=0.69U NW=0.3U
XI10 NET80 NET55 IVG PW=0.84U NW=0.56U
.ENDS FFSDSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSRHD1X                                                           *
* LAST TIME SAVED: DEC  1 14:35:17 2003                                       *
*******************************************************************************
.SUBCKT FFSDSRHD1X Q QN CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.68U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.68U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.18U
MN0 NET55 SN NET180 GND N18 W=0.54U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET180 NET117 GND GND N18 W=0.54U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=1.1U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.1U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.7U PW=0.7U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=1.2U NW=0.8U
XI5 Q NET80 IVG PW=1.2U NW=0.8U
XI13 NET94 NET115 IVG PW=0.6U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSHDLX                                                            *
* LAST TIME SAVED: DEC  1 14:37:17 2003                                       *
*******************************************************************************
.SUBCKT FFSDSHDLX Q QN CK D SN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=0.84U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=0.72U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=0.72U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.5U PW=0.5U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=0.64U NW=0.42U
XI5 Q NET80 IVG PW=0.64U NW=0.42U
XI13 NET94 NET115 IVG PW=0.42U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:37:00 2003                                       *
*******************************************************************************
.SUBCKT FFSDSHD4X Q QN CK D SN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=1.1U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=2.52U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 SN GND GND N18 W=0.8U L=0.18U
MN3 NET73 SN GND GND N18 W=2.16U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=2.16U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG_1 NW=0.9U PW=1.5U PL0=0.19U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.35U PW=1.35U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.7U PW=0.7U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.8U
XI12 QN NET55 IVG PW=4.8U NW=3.2U
XI5 Q NET80 IVG PW=4.8U NW=3.2U
XI13 NET94 NET115 IVG PW=0.93U NW=0.3U
XI10 NET80 NET55 IVG PW=1.77U NW=1.18U
.ENDS FFSDSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSHD2X                                                            *
* LAST TIME SAVED: DEC 27 18:43:20 2003                                       *
*******************************************************************************
.SUBCKT FFSDSHD2X Q QN CK D SN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=1.72U L=0.19U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=1.57U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.57U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.1U PW=1.1U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.45U
XI12 QN NET55 IVG PW=2.4U NW=1.6U
XI5 Q NET80 IVG PW=2.4U NW=1.6U
XI13 NET94 NET115 IVG PW=0.69U NW=0.3U
XI10 NET80 NET55 IVG PW=0.84U NW=0.56U
.ENDS FFSDSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDSHD1X                                                            *
* LAST TIME SAVED: DEC 27 23:23:52 2003                                       *
*******************************************************************************
.SUBCKT FFSDSHD1X Q QN CK D SN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=1.28U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 SN GND GND N18 W=0.6U L=0.18U
MN3 NET73 SN GND GND N18 W=1.1U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.1U L=0.19U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.7U PW=0.7U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=1.2U NW=0.8U
XI5 Q NET80 IVG PW=1.2U NW=0.8U
XI13 NET94 NET115 IVG PW=0.6U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDRHDLX                                                            *
* LAST TIME SAVED: DEC 27 23:26:09 2003                                       *
*******************************************************************************
.SUBCKT FFSDRHDLX Q QN CK D RN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.1U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.1U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.19U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 GND GND N18 W=0.3U L=0.18U
MN6 NET55 NET117 GND GND N18 W=0.42U L=0.18U
MN2 NET70 NET96 GND GND N18 W=0.56U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.5U PW=0.5U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=0.64U NW=0.42U
XI5 Q NET80 IVG PW=0.64U NW=0.42U
XI13 NET94 NET115 IVG PW=0.42U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDRHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:38:09 2003                                       *
*******************************************************************************
.SUBCKT FFSDRHD4X Q QN CK D RN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=3.3U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=3.3U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1.68U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 GND GND N18 W=0.3U L=0.18U
MN6 NET55 NET117 GND GND N18 W=0.72U L=0.18U
MN2 NET70 NET96 GND GND N18 W=1.68U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG_1 NW=0.9U PW=1.5U PL0=0.19U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.35U PW=1.35U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.7U PW=0.7U
XI21 NET117 RN IVG PW=1.5U NW=1U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.8U
XI12 QN NET55 IVG PW=4.8U NW=3.2U
XI5 Q NET80 IVG PW=4.8U NW=3.2U
XI13 NET94 NET115 IVG PW=0.93U NW=0.3U
XI10 NET80 NET55 IVG PW=1.77U NW=1.18U
.ENDS FFSDRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDRHD2X                                                            *
* LAST TIME SAVED: DEC  1 14:37:54 2003                                       *
*******************************************************************************
.SUBCKT FFSDRHD2X Q QN CK D RN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=2.25U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=2.25U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=0.86U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 GND GND N18 W=0.3U L=0.18U
MN6 NET55 NET117 GND GND N18 W=0.42U L=0.18U
MN2 NET70 NET96 GND GND N18 W=1.22U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.1U PW=1.1U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.81U NW=0.54U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.45U
XI12 QN NET55 IVG PW=2.4U NW=1.6U
XI5 Q NET80 IVG PW=2.4U NW=1.6U
XI13 NET94 NET115 IVG PW=0.69U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDRHD1X                                                            *
* LAST TIME SAVED: DEC 27 23:25:47 2003                                       *
*******************************************************************************
.SUBCKT FFSDRHD1X Q QN CK D RN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.68U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.68U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.19U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 GND GND N18 W=0.3U L=0.18U
MN6 NET55 NET117 GND GND N18 W=0.42U L=0.18U
MN2 NET70 NET96 GND GND N18 W=0.86U L=0.18U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI36 NET61 D NET76 TE TRIIVG NW=0.54U PW=0.9U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.7U PW=0.7U
XI6 NET61 NET96 NET115 NET94 TG1G NW=0.42U PW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 QN NET55 IVG PW=1.2U NW=0.8U
XI5 Q NET80 IVG PW=1.2U NW=0.8U
XI13 NET94 NET115 IVG PW=0.6U NW=0.3U
XI10 NET80 NET55 IVG PW=0.64U NW=0.42U
.ENDS FFSDRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSRHDLX                                                          *
* LAST TIME SAVED: DEC  1 14:40:31 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSRHDLX Q CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET92 VDD P18 W=0.45U L=0.18U
MP3 NET55 NET117 NET92 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.84U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.1U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.1U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.18U
MN1 NET92 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET92 NET117 GND GND N18 W=0.42U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=0.72U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=0.72U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.32U PW=0.48U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.45U PW=0.51U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET92 NET94 NET115 TG1G NW=0.5U PW=0.5U
XI21 NET117 SN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 Q NET92 IVG PW=0.64U NW=0.42U
XI13 NET94 NET115 IVG PW=0.42U NW=0.3U
XI10 NET80 NET92 IVG PW=0.42U NW=0.3U
.ENDS FFSDQSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSRHD4X                                                          *
* LAST TIME SAVED: DEC  1 14:40:07 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSRHD4X Q CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET92 VDD P18 W=0.45U L=0.18U
MP3 NET55 NET117 NET92 VDD P18 W=1.44U L=0.18U
MP8 VDD RN NET55 VDD P18 W=1.44U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=3.68U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=3.68U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1.68U L=0.18U
MN1 NET92 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET92 NET117 GND GND N18 W=0.72U L=0.18U
MN5 NET142 RN GND GND N18 W=0.8U L=0.18U
MN3 NET73 RN GND GND N18 W=2.32U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=2.32U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.6U PW=0.9U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=1U PW=1.17U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET92 NET94 NET115 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI21 NET117 SN IVG PW=1.5U NW=1U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.75U
XI12 Q NET92 IVG PW=4.8U NW=3.2U
XI13 NET94 NET115 IVG PW=0.9U NW=0.3U
XI10 NET80 NET92 IVG PW=0.42U NW=0.3U
.ENDS FFSDQSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSRHD2X                                                          *
* LAST TIME SAVED: DEC  1 14:39:36 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSRHD2X Q CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET92 VDD P18 W=0.45U L=0.18U
MP3 NET55 NET117 NET92 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.84U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=2.25U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=2.25U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=0.86U L=0.18U
MN1 NET92 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET92 NET117 GND GND N18 W=0.42U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=1.57U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.57U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.42U PW=0.64U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.51U PW=0.69U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET92 NET94 NET115 TG1G NW=1.1U PW=1.1U
XI21 NET117 SN IVG PW=0.81U NW=0.54U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.45U
XI12 Q NET92 IVG PW=2.4U NW=1.6U
XI13 NET94 NET115 IVG PW=0.69U NW=0.3U
XI10 NET80 NET92 IVG PW=0.42U NW=0.3U
.ENDS FFSDQSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSRHD1X                                                          *
* LAST TIME SAVED: DEC  1 14:39:11 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSRHD1X Q CK D RN SN TE TI
MP5 NET143 NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET92 VDD P18 W=0.45U L=0.18U
MP3 NET55 NET117 NET92 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.84U L=0.18U
MP6 NET49 NET96 NET70 VDD P18 W=1.68U L=0.18U
MP1 VDD NET117 NET49 VDD P18 W=1.68U L=0.18U
MP7 VDD NET117 NET143 VDD P18 W=1U L=0.18U
MN1 NET92 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN6 NET92 NET117 GND GND N18 W=0.42U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=1.1U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.1U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.42U PW=0.64U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.42U PW=0.64U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET92 NET94 NET115 TG1G NW=0.7U PW=0.7U
XI21 NET117 SN IVG PW=0.64U NW=0.42U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 Q NET92 IVG PW=1.2U NW=0.8U
XI13 NET94 NET115 IVG PW=0.6U NW=0.3U
XI10 NET80 NET92 IVG PW=0.42U NW=0.3U
.ENDS FFSDQSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSHDLX                                                           *
* LAST TIME SAVED: DEC  1 14:42:36 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSHDLX Q CK D SN TE TI
XI34 NET81 NET54 NET98 NET79 TRIIVG NW=0.45U PW=0.51U
XI31 NET81 NET46 NET79 NET98 TRIIVG NW=0.3U PW=0.42U
XI33 NET54 TI TE NET69 TRIIVG NW=0.3U PW=0.42U
XI32 NET54 D NET69 TE TRIIVG NW=0.32U PW=0.48U
MP1 VDD NET102 NET59 VDD P18 W=1.1U L=0.18U
MP5 VDD NET102 NET53 VDD P18 W=1U L=0.18U
MP7 NET53 NET66 NET50 VDD P18 W=0.6U L=0.18U
MP6 NET59 NET81 NET46 VDD P18 W=1.1U L=0.18U
MP4 NET50 NET79 NET77 VDD P18 W=0.6U L=0.18U
MN5 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET77 NET98 NET68 GND N18 W=0.3U L=0.18U
MN3 NET46 NET81 GND GND N18 W=0.56U L=0.18U
MN6 NET77 NET102 GND GND N18 W=0.42U L=0.18U
XI9 NET46 NET77 NET79 NET98 TG1G NW=0.5U PW=0.5U
XI12 Q NET77 IVG PW=0.64U NW=0.42U
XI10 NET66 NET77 IVG PW=0.42U NW=0.3U
XI21 NET102 SN IVG PW=0.64U NW=0.42U
XI13 NET79 NET98 IVG PW=0.42U NW=0.3U
XI4 NET98 CK IVG PW=0.3U NW=0.3U
XI20 NET69 TE IVG PW=0.42U NW=0.3U
.ENDS FFSDQSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:42:14 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSHD4X Q CK D SN TE TI
XI34 NET81 NET54 NET98 NET79 TRIIVG NW=1U PW=1.17U
XI31 NET81 NET46 NET79 NET98 TRIIVG NW=0.3U PW=0.42U
XI33 NET54 TI TE NET69 TRIIVG NW=0.3U PW=0.42U
XI32 NET54 D NET69 TE TRIIVG NW=0.6U PW=0.9U
MP1 VDD NET102 NET59 VDD P18 W=3.68U L=0.18U
MP5 VDD NET102 NET53 VDD P18 W=1.68U L=0.18U
MP7 NET53 NET66 NET50 VDD P18 W=0.6U L=0.18U
MP6 NET59 NET81 NET46 VDD P18 W=3.68U L=0.18U
MP4 NET50 NET79 NET77 VDD P18 W=0.6U L=0.18U
MN5 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET77 NET98 NET68 GND N18 W=0.3U L=0.18U
MN3 NET46 NET81 GND GND N18 W=1.81U L=0.18U
MN6 NET77 NET102 GND GND N18 W=0.72U L=0.18U
XI9 NET46 NET77 NET79 NET98 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI12 Q NET77 IVG PW=4.8U NW=3.2U
XI10 NET66 NET77 IVG PW=0.42U NW=0.3U
XI21 NET102 SN IVG PW=1.5U NW=1U
XI13 NET79 NET98 IVG PW=0.9U NW=0.3U
XI4 NET98 CK IVG PW=0.3U NW=0.75U
XI20 NET69 TE IVG PW=0.42U NW=0.3U
.ENDS FFSDQSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSHD2X                                                           *
* LAST TIME SAVED: DEC  1 14:41:48 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSHD2X Q CK D SN TE TI
XI34 NET81 NET54 NET98 NET79 TRIIVG NW=0.51U PW=0.96U
XI31 NET81 NET46 NET79 NET98 TRIIVG NW=0.3U PW=0.42U
XI33 NET54 TI TE NET69 TRIIVG NW=0.3U PW=0.42U
XI32 NET54 D NET69 TE TRIIVG NW=0.42U PW=0.64U
MP1 VDD NET102 NET59 VDD P18 W=2.25U L=0.18U
MP5 VDD NET102 NET53 VDD P18 W=0.86U L=0.18U
MP7 NET53 NET66 NET50 VDD P18 W=0.6U L=0.18U
MP6 NET59 NET81 NET46 VDD P18 W=2.25U L=0.18U
MP4 NET50 NET79 NET77 VDD P18 W=0.6U L=0.18U
MN5 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET77 NET98 NET68 GND N18 W=0.3U L=0.18U
MN3 NET46 NET81 GND GND N18 W=1.22U L=0.18U
MN6 NET77 NET102 GND GND N18 W=0.42U L=0.18U
XI9 NET46 NET77 NET79 NET98 TG1G NW=1.1U PW=1.1U
XI12 Q NET77 IVG PW=2.4U NW=1.6U
XI10 NET66 NET77 IVG PW=0.42U NW=0.3U
XI21 NET102 SN IVG PW=0.81U NW=0.54U
XI13 NET79 NET98 IVG PW=0.69U NW=0.3U
XI4 NET98 CK IVG PW=0.3U NW=0.45U
XI20 NET69 TE IVG PW=0.42U NW=0.3U
.ENDS FFSDQSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQSHD1X                                                           *
* LAST TIME SAVED: DEC  1 14:41:23 2003                                       *
*******************************************************************************
.SUBCKT FFSDQSHD1X Q CK D SN TE TI
XI34 NET81 NET54 NET98 NET79 TRIIVG NW=0.42U PW=0.64U
XI31 NET81 NET46 NET79 NET98 TRIIVG NW=0.3U PW=0.42U
XI33 NET54 TI TE NET69 TRIIVG NW=0.3U PW=0.42U
XI32 NET54 D NET69 TE TRIIVG NW=0.42U PW=0.64U
MP1 VDD NET102 NET59 VDD P18 W=1.68U L=0.18U
MP5 VDD NET102 NET53 VDD P18 W=1U L=0.18U
MP7 NET53 NET66 NET50 VDD P18 W=0.6U L=0.18U
MP6 NET59 NET81 NET46 VDD P18 W=1.68U L=0.18U
MP4 NET50 NET79 NET77 VDD P18 W=0.6U L=0.18U
MN5 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET77 NET98 NET68 GND N18 W=0.3U L=0.18U
MN3 NET46 NET81 GND GND N18 W=0.86U L=0.18U
MN6 NET77 NET102 GND GND N18 W=0.42U L=0.18U
XI9 NET46 NET77 NET79 NET98 TG1G NW=0.7U PW=0.7U
XI12 Q NET77 IVG PW=1.2U NW=0.8U
XI10 NET66 NET77 IVG PW=0.42U NW=0.3U
XI21 NET102 SN IVG PW=0.64U NW=0.42U
XI13 NET79 NET98 IVG PW=0.6U NW=0.3U
XI4 NET98 CK IVG PW=0.3U NW=0.3U
XI20 NET69 TE IVG PW=0.42U NW=0.3U
.ENDS FFSDQSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQRHDLX                                                           *
* LAST TIME SAVED: DEC  1 14:44:27 2003                                       *
*******************************************************************************
.SUBCKT FFSDQRHDLX Q CK D RN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=0.84U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=0.72U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=0.72U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.32U PW=0.48U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.45U PW=0.51U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.5U PW=0.5U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 Q NET55 IVG PW=0.64U NW=0.42U
XI13 NET94 NET115 IVG PW=0.42U NW=0.3U
XI10 NET80 NET55 IVG PW=0.42U NW=0.3U
.ENDS FFSDQRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQRHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:43:58 2003                                       *
*******************************************************************************
.SUBCKT FFSDQRHD4X Q CK D RN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET55 VDD P18 W=1.1U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=2.81U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 RN GND GND N18 W=0.8U L=0.18U
MN3 NET73 RN GND GND N18 W=2.32U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=2.32U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.6U PW=0.9U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=1U PW=1.17U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.75U
XI12 Q NET55 IVG PW=4.8U NW=3.2U
XI13 NET94 NET115 IVG PW=0.9U NW=0.3U
XI10 NET80 NET55 IVG PW=0.42U NW=0.3U
.ENDS FFSDQRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQRHD2X                                                           *
* LAST TIME SAVED: DEC  1 14:43:32 2003                                       *
*******************************************************************************
.SUBCKT FFSDQRHD2X Q CK D RN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=1.72U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=1.57U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.57U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.42U PW=0.64U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.51U PW=0.69U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET55 NET94 NET115 TG1G NW=1.1U PW=1.1U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.45U
XI12 Q NET55 IVG PW=2.4U NW=1.6U
XI13 NET94 NET115 IVG PW=0.69U NW=0.3U
XI10 NET80 NET55 IVG PW=0.42U NW=0.3U
.ENDS FFSDQRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQRHD1X                                                           *
* LAST TIME SAVED: DEC  1 14:43:08 2003                                       *
*******************************************************************************
.SUBCKT FFSDQRHD1X Q CK D RN TE TI
MP5 VDD NET80 NET58 VDD P18 W=0.45U L=0.18U
MP4 NET58 NET94 NET55 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET55 VDD P18 W=0.64U L=0.18U
MP6 VDD NET96 NET70 VDD P18 W=1.28U L=0.18U
MN1 NET55 NET115 NET82 GND N18 W=0.3U L=0.18U
MN4 NET82 NET80 NET142 GND N18 W=0.3U L=0.18U
MN5 NET142 RN GND GND N18 W=0.6U L=0.18U
MN3 NET73 RN GND GND N18 W=1.1U L=0.18U
MN2 NET70 NET96 NET73 GND N18 W=1.1U L=0.18U
XI36 NET61 D NET76 TE TRIIVG NW=0.42U PW=0.64U
XI33 NET96 NET70 NET94 NET115 TRIIVG NW=0.3U PW=0.42U
XI38 NET96 NET61 NET115 NET94 TRIIVG NW=0.42U PW=0.64U
XI37 NET61 TI TE NET76 TRIIVG NW=0.3U PW=0.42U
XI9 NET70 NET55 NET94 NET115 TG1G NW=0.7U PW=0.7U
XI20 NET76 TE IVG PW=0.42U NW=0.3U
XI4 NET115 CK IVG PW=0.3U NW=0.3U
XI12 Q NET55 IVG PW=1.2U NW=0.8U
XI13 NET94 NET115 IVG PW=0.6U NW=0.3U
XI10 NET80 NET55 IVG PW=0.42U NW=0.3U
.ENDS FFSDQRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQHDLX                                                            *
* LAST TIME SAVED: DEC  1 14:45:43 2003                                       *
*******************************************************************************
.SUBCKT FFSDQHDLX Q CK D TE TI
XI21 NET33 NET43 NET32 NET24 TRIIVG NW=0.45U PW=0.51U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET43 D NET57 TE TRIIVG NW=0.32U PW=0.48U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET43 TI TE NET57 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI20 NET57 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSDQHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:45:18 2003                                       *
*******************************************************************************
.SUBCKT FFSDQHD4X Q CK D TE TI
XI21 NET33 NET43 NET32 NET24 TRIIVG NW=1U PW=1.17U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET43 D NET57 TE TRIIVG NW=0.6U PW=0.9U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET43 TI TE NET57 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI20 NET57 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.81U NW=1.81U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
.ENDS FFSDQHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQHD2X                                                            *
* LAST TIME SAVED: DEC  1 14:45:02 2003                                       *
*******************************************************************************
.SUBCKT FFSDQHD2X Q CK D TE TI
XI21 NET33 NET43 NET32 NET24 TRIIVG NW=0.51U PW=0.69U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET43 D NET57 TE TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET43 TI TE NET57 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI20 NET57 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFSDQHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDQHD1X                                                            *
* LAST TIME SAVED: DEC  1 14:44:46 2003                                       *
*******************************************************************************
.SUBCKT FFSDQHD1X Q CK D TE TI
XI21 NET33 NET43 NET32 NET24 TRIIVG NW=0.42U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET43 D NET57 TE TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET43 TI TE NET57 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI20 NET57 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSDQHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSRHDLX                                                          *
* LAST TIME SAVED: DEC  1 14:47:07 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSRHDLX Q QN CKN D RN SN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=1.01U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=1.01U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=0.81U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.58U L=0.18U
MN6 NET53 SN NET191 GND N18 W=0.58U L=0.18U
MN3 NET83 SN GND GND N18 W=0.81U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET53 NET92 NET93 TG1G NW=0.5U PW=0.5U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=0.64U NW=0.42U
XI4 NET92 CKN IVG PW=0.9U NW=0.3U
XI5 Q NET66 IVG PW=0.64U NW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI10 NET66 NET53 IVG PW=0.42U NW=0.3U
.ENDS FFSDNSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSRHD4X                                                          *
* LAST TIME SAVED: DEC 27 23:16:58 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSRHD4X Q QN CKN D RN SN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=1.1U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=2.82U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=2.82U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1.68U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.8U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=2.25U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.92U L=0.18U
MN6 NET53 SN NET191 GND N18 W=0.92U L=0.18U
MN3 NET83 SN GND GND N18 W=2.25U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.45U PW=1.62U
XI9 NET80 NET53 NET92 NET93 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.7U PW=0.7U
XI13 NET93 NET92 IVG PW=0.3U NW=0.48U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=4.8U NW=3.2U
XI4 NET92 CKN IVG PW=1.44U NW=0.3U
XI5 Q NET66 IVG PW=4.8U NW=3.2U
XI21 NET117 RN IVG PW=1.5U NW=1U
XI10 NET66 NET53 IVG PW=1.77U NW=1.18U
.ENDS FFSDNSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSRHD2X                                                          *
* LAST TIME SAVED: DEC  1 14:46:23 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSRHD2X Q QN CKN D RN SN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=2.04U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=2.04U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=0.86U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=1.74U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.58U L=0.18U
MN6 NET53 SN NET191 GND N18 W=0.58U L=0.18U
MN3 NET83 SN GND GND N18 W=1.74U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=1.05U
XI9 NET80 NET53 NET92 NET93 TG1G NW=1.1U PW=1.1U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.5U PW=0.5U
XI13 NET93 NET92 IVG PW=0.3U NW=0.45U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=2.4U NW=1.6U
XI4 NET92 CKN IVG PW=1.2U NW=0.3U
XI5 Q NET66 IVG PW=2.4U NW=1.6U
XI21 NET117 RN IVG PW=0.81U NW=0.54U
XI10 NET66 NET53 IVG PW=0.84U NW=0.56U
.ENDS FFSDNSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSRHD1X                                                          *
* LAST TIME SAVED: DEC 27 23:07:01 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSRHD1X Q QN CKN D RN SN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=1.56U L=0.19U
MP1 VDD NET117 NET62 VDD P18 W=1.56U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=1.22U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.58U L=0.18U
MN6 NET53 SN NET191 GND N18 W=0.58U L=0.18U
MN3 NET83 SN GND GND N18 W=1.22U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET53 NET92 NET93 TG1G NW=0.7U PW=0.7U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=1.2U NW=0.8U
XI4 NET92 CKN IVG PW=0.78U NW=0.3U
XI5 Q NET66 IVG PW=1.2U NW=0.8U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI10 NET66 NET53 IVG PW=0.64U NW=0.42U
.ENDS FFSDNSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSHDLX                                                           *
* LAST TIME SAVED: DEC  1 14:48:17 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSHDLX Q QN CKN D SN TE TI
MP5 VDD NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 VDD NET94 NET80 VDD P18 W=0.77U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=0.81U L=0.18U
MN3 NET83 SN GND GND N18 W=0.81U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET53 NET92 NET93 TG1G NW=0.5U PW=0.5U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=0.64U NW=0.42U
XI4 NET92 CKN IVG PW=0.9U NW=0.3U
XI5 Q NET66 IVG PW=0.64U NW=0.42U
XI10 NET66 NET53 IVG PW=0.42U NW=0.3U
.ENDS FFSDNSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:48:01 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSHD4X Q QN CKN D SN TE TI
MP5 VDD NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=1.1U L=0.18U
MP6 VDD NET94 NET80 VDD P18 W=2.15U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.8U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=2.25U L=0.18U
MN3 NET83 SN GND GND N18 W=2.25U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG_1 NW=0.45U PW=1.62U PL0=0.19U
XI9 NET80 NET53 NET92 NET93 TG1G NW=1.35U PW=1.35U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.7U PW=0.7U
XI13 NET93 NET92 IVG PW=0.3U NW=0.48U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=4.8U NW=3.2U
XI4 NET92 CKN IVG PW=1.44U NW=0.3U
XI5 Q NET66 IVG PW=4.8U NW=3.2U
XI10 NET66 NET53 IVG PW=1.77U NW=1.18U
.ENDS FFSDNSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSHD2X                                                           *
* LAST TIME SAVED: DEC 27 23:07:27 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSHD2X Q QN CKN D SN TE TI
MP5 VDD NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 VDD NET94 NET80 VDD P18 W=1.55U L=0.19U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=1.74U L=0.18U
MN3 NET83 SN GND GND N18 W=1.74U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=1.05U
XI9 NET80 NET53 NET92 NET93 TG1G NW=1.1U PW=1.1U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.5U PW=0.5U
XI13 NET93 NET92 IVG PW=0.3U NW=0.45U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=2.4U NW=1.6U
XI4 NET92 CKN IVG PW=1.2U NW=0.3U
XI5 Q NET66 IVG PW=2.4U NW=1.6U
XI10 NET66 NET53 IVG PW=0.84U NW=0.56U
.ENDS FFSDNSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNSHD1X                                                           *
* LAST TIME SAVED: DEC  1 14:47:30 2003                                       *
*******************************************************************************
.SUBCKT FFSDNSHD1X Q QN CKN D SN TE TI
MP5 VDD NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET53 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET53 VDD P18 W=0.64U L=0.18U
MP6 VDD NET94 NET80 VDD P18 W=1.19U L=0.18U
MN4 NET68 NET66 NET71 GND N18 W=0.3U L=0.18U
MN5 NET71 SN GND GND N18 W=0.6U L=0.18U
MN1 NET53 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 NET83 GND N18 W=1.22U L=0.18U
MN3 NET83 SN GND GND N18 W=1.22U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET53 NET92 NET93 TG1G NW=0.7U PW=0.7U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET53 IVG PW=1.2U NW=0.8U
XI4 NET92 CKN IVG PW=0.78U NW=0.3U
XI5 Q NET66 IVG PW=1.2U NW=0.8U
XI10 NET66 NET53 IVG PW=0.64U NW=0.42U
.ENDS FFSDNSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNRHDLX                                                           *
* LAST TIME SAVED: DEC 27 23:25:24 2003                                       *
*******************************************************************************
.SUBCKT FFSDNRHDLX Q QN CKN D RN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET191 VDD P18 W=0.45U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=1.01U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=1.01U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1U L=0.19U
MN4 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET191 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 GND GND N18 W=0.63U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.42U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET191 NET92 NET93 TG1G NW=0.5U PW=0.5U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET191 IVG PW=0.64U NW=0.42U
XI4 NET92 CKN IVG PW=0.9U NW=0.3U
XI5 Q NET66 IVG PW=0.64U NW=0.42U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI10 NET66 NET191 IVG PW=0.42U NW=0.3U
.ENDS FFSDNRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNRHD4X                                                           *
* LAST TIME SAVED: DEC  1 14:49:05 2003                                       *
*******************************************************************************
.SUBCKT FFSDNRHD4X Q QN CKN D RN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET191 VDD P18 W=0.45U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=2.82U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=2.82U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1.68U L=0.18U
MN4 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET191 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 GND GND N18 W=1.75U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.72U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG_1 NW=0.45U PW=1.62U PL0=0.19U
XI9 NET80 NET191 NET92 NET93 TG1G NW=1.35U PW=1.35U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.7U PW=0.7U
XI13 NET93 NET92 IVG PW=0.3U NW=0.48U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET191 IVG PW=4.8U NW=3.2U
XI4 NET92 CKN IVG PW=1.44U NW=0.3U
XI5 Q NET66 IVG PW=4.8U NW=3.2U
XI21 NET117 RN IVG PW=1.5U NW=1U
XI10 NET66 NET191 IVG PW=1.77U NW=1.18U
.ENDS FFSDNRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNRHD2X                                                           *
* LAST TIME SAVED: DEC  1 14:48:49 2003                                       *
*******************************************************************************
.SUBCKT FFSDNRHD2X Q QN CKN D RN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET191 VDD P18 W=0.45U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=2.04U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=2.04U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=0.86U L=0.18U
MN4 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET191 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 GND GND N18 W=1.35U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.42U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=1.05U
XI9 NET80 NET191 NET92 NET93 TG1G NW=1.1U PW=1.1U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.5U PW=0.5U
XI13 NET93 NET92 IVG PW=0.3U NW=0.45U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET191 IVG PW=2.4U NW=1.6U
XI4 NET92 CKN IVG PW=1.2U NW=0.3U
XI5 Q NET66 IVG PW=2.4U NW=1.6U
XI21 NET117 RN IVG PW=0.81U NW=0.54U
XI10 NET66 NET191 IVG PW=0.84U NW=0.56U
.ENDS FFSDNRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNRHD1X                                                           *
* LAST TIME SAVED: DEC 27 23:25:00 2003                                       *
*******************************************************************************
.SUBCKT FFSDNRHD1X Q QN CKN D RN TE TI
MP5 NET47 NET66 NET50 VDD P18 W=0.45U L=0.18U
MP4 NET50 NET92 NET191 VDD P18 W=0.45U L=0.18U
MP6 NET62 NET94 NET80 VDD P18 W=1.56U L=0.18U
MP1 VDD NET117 NET62 VDD P18 W=1.56U L=0.18U
MP7 VDD NET117 NET47 VDD P18 W=1U L=0.19U
MN4 NET68 NET66 GND GND N18 W=0.3U L=0.18U
MN1 NET191 NET93 NET68 GND N18 W=0.3U L=0.18U
MN2 NET80 NET94 GND GND N18 W=0.95U L=0.18U
MN0 NET191 NET117 GND GND N18 W=0.42U L=0.18U
XI33 NET94 NET80 NET92 NET93 TRIIVG NW=0.3U PW=0.42U
XI37 NET60 TI TE NET75 TRIIVG NW=0.3U PW=0.42U
XI36 NET60 D NET75 TE TRIIVG NW=0.3U PW=0.9U
XI9 NET80 NET191 NET92 NET93 TG1G NW=0.7U PW=0.7U
XI6 NET60 NET94 NET93 NET92 TG1G NW=0.42U PW=0.42U
XI13 NET93 NET92 IVG PW=0.3U NW=0.3U
XI20 NET75 TE IVG PW=0.42U NW=0.3U
XI12 QN NET191 IVG PW=1.2U NW=0.8U
XI4 NET92 CKN IVG PW=0.78U NW=0.3U
XI5 Q NET66 IVG PW=1.2U NW=0.8U
XI21 NET117 RN IVG PW=0.64U NW=0.42U
XI10 NET66 NET191 IVG PW=0.64U NW=0.42U
.ENDS FFSDNRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNHDLX                                                            *
* LAST TIME SAVED: DEC  1 14:50:27 2003                                       *
*******************************************************************************
.SUBCKT FFSDNHDLX Q QN CKN D TE TI
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET44 TI TE NET59 TRIIVG NW=0.3U PW=0.42U
XI18 NET44 D NET59 TE TRIIVG NW=0.3U PW=0.9U
XI6 NET44 NET33 NET24 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=0.5U PW=0.5U
XI20 NET59 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.77U NW=0.63U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 CKN IVG PW=0.9U NW=0.3U
.ENDS FFSDNHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:50:11 2003                                       *
*******************************************************************************
.SUBCKT FFSDNHD4X Q QN CKN D TE TI
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET44 TI TE NET59 TRIIVG NW=0.3U PW=0.42U
XI18 NET44 D NET59 TE TRIIVG NW=0.45U PW=1.62U
XI6 NET44 NET33 NET24 NET32 TG1G NW=0.7U PW=0.7U
XI9 NET46 NETQ NET32 NET24 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI20 NET59 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.15U NW=1.75U
XI13 NET24 NET32 IVG PW=0.3U NW=0.48U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CKN IVG PW=1.44U NW=0.3U
.ENDS FFSDNHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNHD2X                                                            *
* LAST TIME SAVED: DEC  1 14:49:56 2003                                       *
*******************************************************************************
.SUBCKT FFSDNHD2X Q QN CKN D TE TI
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET44 TI TE NET59 TRIIVG NW=0.3U PW=0.42U
XI18 NET44 D NET59 TE TRIIVG NW=0.3U PW=1.05U
XI6 NET44 NET33 NET24 NET32 TG1G NW=0.5U PW=0.5U
XI9 NET46 NETQ NET32 NET24 TG1G NW=1.1U PW=1.1U
XI20 NET59 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.55U NW=1.35U PL=0.18U NL=0.19U
XI13 NET24 NET32 IVG PW=0.3U NW=0.45U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CKN IVG PW=1.2U NW=0.3U
.ENDS FFSDNHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDNHD1X                                                            *
* LAST TIME SAVED: DEC  1 14:49:41 2003                                       *
*******************************************************************************
.SUBCKT FFSDNHD1X Q QN CKN D TE TI
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET44 TI TE NET59 TRIIVG NW=0.3U PW=0.42U
XI18 NET44 D NET59 TE TRIIVG NW=0.3U PW=0.9U
XI6 NET44 NET33 NET24 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=0.7U PW=0.7U
XI20 NET59 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.19U NW=0.95U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CKN IVG PW=0.78U NW=0.3U
.ENDS FFSDNHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDHDLX                                                             *
* LAST TIME SAVED: NOV 21 10:51:57 2003                                       *
*******************************************************************************
.SUBCKT FFSDHDLX Q QN CK D TE TI
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET47 TI TE NET62 TRIIVG NW=0.3U PW=0.42U
XI18 NET47 D NET62 TE TRIIVG NW=0.54U PW=0.9U
XI6 NET47 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI20 NET62 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.54U NW=0.36U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSDHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDHD4X                                                             *
* LAST TIME SAVED: NOV 21 10:04:56 2003                                       *
*******************************************************************************
.SUBCKT FFSDHD4X Q QN CK D TE TI
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET47 TI TE NET62 TRIIVG NW=0.3U PW=0.42U
XI18 NET47 D NET62 TE TRIIVG_1 NW=0.9U PW=1.5U PL0=0.19U
XI6 NET47 NET33 NET32 NET24 TG1G NW=0.7U PW=0.7U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI20 NET62 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.52U NW=1.68U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
.ENDS FFSDHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDHD2XSPG                                                          *
* LAST TIME SAVED: NOV 21 09:46:39 2003                                       *
*******************************************************************************
.SUBCKT FFSDHD2XSPG Q QN CK D TE TI
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET47 TI TE NET62 TRIIVG NW=0.3U PW=0.42U
XI18 NET47 D NET62 TE TRIIVG NW=0.54U PW=0.9U
XI6 NET47 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI20 NET62 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFSDHD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDHD2X                                                             *
* LAST TIME SAVED: NOV 20 19:30:32 2003                                       *
*******************************************************************************
.SUBCKT FFSDHD2X Q QN CK D TE TI
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET47 TI TE NET62 TRIIVG NW=0.3U PW=0.42U
XI18 NET47 D NET62 TE TRIIVG NW=0.54U PW=0.9U
XI6 NET47 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI20 NET62 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFSDHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDHD1X                                                             *
* LAST TIME SAVED: NOV 20 17:22:25 2003                                       *
*******************************************************************************
.SUBCKT FFSDHD1X Q QN CK D TE TI
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI19 NET47 TI TE NET62 TRIIVG NW=0.3U PW=0.42U
XI18 NET47 D NET62 TE TRIIVG NW=0.54U PW=0.9U
XI6 NET47 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI20 NET62 TE IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFSDHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDCRHDLX                                                           *
* LAST TIME SAVED: MAR  4 15:10:51 2003                                       *
*******************************************************************************
.SUBCKT FFSDCRHDLX Q QN CK D RN TE TI
XI18 NET63 RN D ND2G PW=0.6U NW=0.5U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI25 NET72 NET51 TE NET68 TG1G NW=0.42U PW=0.42U
XI6 NET51 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI19 NET63 NET51 NET68 TE TG1G NW=0.8U PW=0.8U
XI21 NET72 TI IVG PW=0.42U NW=0.3U
XI20 NET68 TE IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=0.64U NW=0.42U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFSDCRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDCRHD4X                                                           *
* LAST TIME SAVED: MAR  4 15:10:33 2003                                       *
*******************************************************************************
.SUBCKT FFSDCRHD4X Q QN CK D RN TE TI
XI18 NET63 RN D ND2G PW=1.47U NW=1.18U
XI17 NET33 NET46 NET32 NET122 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET122 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET63 NET51 NET66 TE TG1G NW=0.8U PW=0.8U
XI25 NET74 NET51 TE NET66 TG1G NW=0.42U PW=0.42U
XI6 NET51 NET33 NET122 NET32 TG1G NW=0.8U PW=0.8U
XI9 NET46 NETQN NET32 NET122 TG1G NW=1.18U PW=1.18U
XI7 NET46 NET33 IVG PW=3.44U NW=2.3U
XI20 NET66 TE IVG PW=0.64U NW=0.42U
XI13 NET32 NET122 IVG PW=0.96U NW=0.48U
XI12 QN NETQN IVG PW=4.8U NW=3.2U
XI10 NETQ NETQN IVG PW=1.68U NW=1.14U
XI21 NET74 TI IVG PW=0.42U NW=0.3U
XI5 Q NETQ IVG PW=4.8U NW=3.2U
XI4 NET122 CK IVG PW=1.2U NW=0.6U
.ENDS FFSDCRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDCRHD2X                                                           *
* LAST TIME SAVED: MAR  4 15:10:14 2003                                       *
*******************************************************************************
.SUBCKT FFSDCRHD2X Q QN CK D RN TE TI
XI18 NET63 RN D ND2G PW=0.96U NW=0.8U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET63 NET51 NET66 TE TG1G NW=0.8U PW=0.8U
XI25 NET73 NET51 TE NET66 TG1G NW=0.42U PW=0.42U
XI6 NET51 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI21 NET73 TI IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI20 NET66 TE IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFSDCRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFSDCRHD1X                                                           *
* LAST TIME SAVED: MAR  4 15:09:57 2003                                       *
*******************************************************************************
.SUBCKT FFSDCRHD1X Q QN CK D RN TE TI
XI18 NET34 RN D ND2G PW=0.66U NW=0.55U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET53 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI25 NET120 NET53 TE NET70 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI19 NET34 NET53 NET70 TE TG1G NW=0.8U PW=0.8U
XI21 NET120 TI IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI20 NET70 TE IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=1.2U NW=0.8U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFSDCRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSRHDLX                                                           *
* LAST TIME SAVED: MAR 13 15:07:12 2003                                       *
*******************************************************************************
.SUBCKT FFJKSRHDLX Q QN CK J K RN SN
XI21 NET66 SN IVG PW=0.64U NW=0.42U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET112 NETQ IVG PW=0.64U NW=0.42U
XI5 QN NET112 IVG PW=0.64U NW=0.42U
XI13 NET67 NET164 IVG PW=0.6U NW=0.3U
XI4 NET164 CK IVG PW=0.84U NW=0.42U
XI9 NET120 NETQ NET67 NET164 TG1G NW=0.7U PW=0.7U
XI6 NET39 NET69 NET164 NET67 TG1G NW=0.42U PW=0.42U
XI33 NET69 NET120 NET67 NET164 TRIIVG NW=0.3U PW=0.42U
MP0 NET99 NET67 NETQ VDD P18 W=0.45U L=0.18U
MP1 NET84 NET66 NETQ VDD P18 W=0.84U L=0.18U
MP2 VDD NET66 NET87 VDD P18 W=1.16U L=0.18U
MP8 VDD RN NET84 VDD P18 W=0.84U L=0.18U
MP6 NET93 NET112 NET99 VDD P18 W=0.45U L=0.18U
MP7 VDD NET66 NET93 VDD P18 W=1U L=0.18U
MP9 NET87 NET69 NET120 VDD P18 W=1.16U L=0.18U
MP4 NET40 NETQ NET39 VDD P18 W=1.2U L=0.18U
MP5 VDD NET62 NET39 VDD P18 W=0.72U L=0.18U
MP3 VDD K NET40 VDD P18 W=1.2U L=0.18U
MN5 NET126 RN GND GND N18 W=0.6U L=0.18U
MN6 NETQ NET66 GND GND N18 W=0.42U L=0.18U
MN0 NET123 RN GND GND N18 W=0.77U L=0.18U
MN4 NET120 NET69 NET123 GND N18 W=0.77U L=0.18U
MN7 NETQ NET164 NET114 GND N18 W=0.3U L=0.18U
MN8 NET114 NET112 NET126 GND N18 W=0.3U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.6U L=0.18U
MN2 NET52 K GND GND N18 W=0.6U L=0.18U
MN1 NET39 NET62 NET52 GND N18 W=0.6U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSRHD4X                                                           *
* LAST TIME SAVED: MAR 13 14:45:55 2003                                       *
*******************************************************************************
.SUBCKT FFJKSRHD4X Q QN CK J K RN SN
XI21 NET174 SN IVG PW=1.5U NW=1U
XI12 Q NET255 IVG PW=4.8U NW=3.2U
XI10 NET242 NET255 IVG PW=1.68U NW=1.14U
XI5 QN NET242 IVG PW=4.8U NW=3.2U
XI13 NET189 NET190 IVG PW=0.96U NW=0.48U
XI4 NET190 CK IVG PW=1.2U NW=0.6U
XI9 NET247 NET255 NET189 NET190 TG1G NW=1.18U PW=1.18U
XI6 NET198 NET191 NET190 NET189 TG1G NW=0.6U PW=0.6U
XI33 NET191 NET247 NET189 NET190 TRIIVG NW=0.3U PW=0.42U
MP4 NET199 NET255 NET198 VDD P18 W=2.4U L=0.18U
MP5 VDD NET256 NET198 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET199 VDD P18 W=2.4U L=0.18U
MP2 VDD NET174 NET223 VDD P18 W=3.3U L=0.18U
MP7 VDD NET174 NET226 VDD P18 W=1.68U L=0.18U
MP9 NET214 NET174 NET255 VDD P18 W=1.44U L=0.18U
MP0 NET217 NET189 NET255 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET214 VDD P18 W=1.44U L=0.18U
MP6 NET223 NET191 NET247 VDD P18 W=3.3U L=0.18U
MP1 NET226 NET242 NET217 VDD P18 W=0.45U L=0.18U
MN2 NET229 K GND GND N18 W=1.18U L=0.18U
MN1 NET198 NET256 NET229 GND N18 W=1.18U L=0.18U
MN3 NET229 NET255 GND GND N18 W=1.18U L=0.18U
MN7 NET238 RN GND GND N18 W=2.3U L=0.18U
MN6 NET255 NET174 GND GND N18 W=0.72U L=0.18U
MN8 NET244 NET242 NET253 GND N18 W=0.3U L=0.18U
MN0 NET247 NET191 NET238 GND N18 W=2.3U L=0.18U
MN4 NET255 NET190 NET244 GND N18 W=0.3U L=0.18U
MN5 NET253 RN GND GND N18 W=0.8U L=0.18U
XI18 NET256 NET255 J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSRHD2X                                                           *
* LAST TIME SAVED: MAR 13 15:03:39 2003                                       *
*******************************************************************************
.SUBCKT FFJKSRHD2X Q QN CK J K RN SN
XI21 NET67 SN IVG PW=0.81U NW=0.54U
XI12 Q NET257 IVG PW=2.4U NW=1.6U
XI10 NET116 NET257 IVG PW=0.84U NW=0.56U
XI5 QN NET116 IVG PW=2.4U NW=1.6U
XI36 NET65 NET63 IVG PW=0.84U NW=0.42U
XI4 NET63 CK IVG PW=1.2U NW=0.6U
XI9 NET121 NET257 NET65 NET63 TG1G NW=1.1U PW=1.1U
XI6 NET45 NET70 NET63 NET65 TG1G NW=0.42U PW=0.42U
XI33 NET70 NET121 NET65 NET63 TRIIVG NW=0.3U PW=0.42U
MP1 NET94 NET116 NET97 VDD P18 W=0.45U L=0.18U
MP2 NET91 NET67 NET257 VDD P18 W=1.2U L=0.18U
MP8 VDD RN NET91 VDD P18 W=1.2U L=0.18U
MP4 NET109 NET257 NET45 VDD P18 W=1.66U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET109 VDD P18 W=1.66U L=0.18U
MP6 NET85 NET70 NET121 VDD P18 W=1.68U L=0.18U
MP9 VDD NET67 NET85 VDD P18 W=1.68U L=0.18U
MP7 VDD NET67 NET94 VDD P18 W=0.86U L=0.18U
MP0 NET97 NET65 NET257 VDD P18 W=0.45U L=0.18U
MN3 NET55 NET257 GND GND N18 W=0.9U L=0.18U
MN4 NET121 NET70 NET124 GND N18 W=1.12U L=0.18U
MN6 NET257 NET67 GND GND N18 W=0.42U L=0.18U
MN5 NET118 NET116 NET115 GND N18 W=0.3U L=0.18U
MN7 NET115 RN GND GND N18 W=0.6U L=0.18U
MN8 NET257 NET63 NET118 GND N18 W=0.3U L=0.18U
MN0 NET124 RN GND GND N18 W=1.12U L=0.18U
MN2 NET55 K GND GND N18 W=0.9U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=0.9U L=0.18U
XI18 NET62 NET257 J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSRHD1X                                                           *
* LAST TIME SAVED: MAR 13 14:36:20 2003                                       *
*******************************************************************************
.SUBCKT FFJKSRHD1X Q QN CK J K RN SN
XI9 NET135 NETQ NET59 NET74 TG1G NW=0.7U PW=0.7U
XI6 NET45 NET61 NET74 NET59 TG1G NW=0.42U PW=0.42U
XI21 NET70 SN IVG PW=0.64U NW=0.42U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NET115 NETQ IVG PW=0.64U NW=0.42U
XI13 NET59 NET74 IVG PW=0.6U NW=0.3U
XI4 NET74 CK IVG PW=0.84U NW=0.42U
XI5 QN NET115 IVG PW=1.2U NW=0.8U
XI34 NET61 NET135 NET59 NET74 TRIIVG NW=0.3U PW=0.42U
MP4 NET107 NETQ NET45 VDD P18 W=1.6U L=0.18U
MP5 VDD NET58 NET45 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET107 VDD P18 W=1.6U L=0.18U
MP1 VDD NET70 NET108 VDD P18 W=1.6U L=0.18U
MP7 VDD NET70 NET90 VDD P18 W=1U L=0.18U
MP0 NET90 NET115 NET87 VDD P18 W=0.45U L=0.18U
MP2 NET87 NET59 NETQ VDD P18 W=0.45U L=0.18U
MP6 NET84 NET70 NETQ VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET84 VDD P18 W=0.84U L=0.18U
MP9 NET108 NET61 NET135 VDD P18 W=1.6U L=0.18U
MN3 NET55 NETQ GND GND N18 W=0.8U L=0.18U
MN0 NETQ NET74 NET117 GND N18 W=0.3U L=0.18U
MN6 NETQ NET70 GND GND N18 W=0.42U L=0.18U
MN2 NET55 K GND GND N18 W=0.8U L=0.18U
MN7 NET129 RN GND GND N18 W=1.06U L=0.18U
MN4 NET117 NET115 NET114 GND N18 W=0.3U L=0.18U
MN1 NET45 NET58 NET55 GND N18 W=0.8U L=0.18U
MN5 NET114 RN GND GND N18 W=0.6U L=0.18U
MN8 NET135 NET61 NET129 GND N18 W=1.06U L=0.18U
XI33 NET58 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSHDLX                                                            *
* LAST TIME SAVED: MAR 13 14:30:28 2003                                       *
*******************************************************************************
.SUBCKT FFJKSHDLX Q QN CK J K SN
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET108 NETQ IVG PW=0.64U NW=0.42U
XI5 QN NET108 IVG PW=0.64U NW=0.42U
XI13 NET66 NET61 IVG PW=0.6U NW=0.3U
XI4 NET61 CK IVG PW=0.84U NW=0.42U
XI21 NET137 SN IVG PW=0.64U NW=0.42U
XI9 NET107 NETQ NET66 NET61 TG1G NW=0.7U PW=0.7U
XI6 NET43 NET68 NET61 NET66 TG1G NW=0.42U PW=0.42U
XI32 NET68 NET107 NET66 NET61 TRIIVG NW=0.3U PW=0.42U
MP4 NET44 NETQ NET43 VDD P18 W=1.2U L=0.18U
MP5 VDD NET65 NET43 VDD P18 W=0.72U L=0.18U
MP3 VDD K NET44 VDD P18 W=1.2U L=0.18U
MP0 NET92 NET66 NETQ VDD P18 W=0.6U L=0.18U
MP1 VDD NET137 NET86 VDD P18 W=1.54U L=0.18U
MP6 NET86 NET68 NET107 VDD P18 W=1.54U L=0.18U
MP7 NET83 NET108 NET92 VDD P18 W=0.6U L=0.18U
MP2 VDD NET137 NET83 VDD P18 W=1U L=0.18U
MN5 NET110 NET108 GND GND N18 W=0.3U L=0.18U
MN3 NET53 NETQ GND GND N18 W=0.6U L=0.18U
MN4 NET107 NET68 GND GND N18 W=0.77U L=0.18U
MN6 NETQ NET137 GND GND N18 W=0.42U L=0.18U
MN0 NETQ NET61 NET110 GND N18 W=0.3U L=0.18U
MN2 NET53 K GND GND N18 W=0.6U L=0.18U
MN1 NET43 NET65 NET53 GND N18 W=0.6U L=0.18U
XI18 NET65 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSHD4X                                                            *
* LAST TIME SAVED: DEC 27 18:42:07 2003                                       *
*******************************************************************************
.SUBCKT FFJKSHD4X Q QN CK J K SN
XI10 NET100 NETQ IVG PW=1.68U NW=1.14U
XI5 QN NET100 IVG PW=4.8U NW=3.2U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI21 NET61 SN IVG PW=1.05U NW=0.7U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
XI32 NET33 NET68 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
MP7 NET72 NET100 NET78 VDD P18 W=0.6U L=0.18U
MP6 NET81 NET33 NET68 VDD P18 W=3.36U L=0.18U
MP2 VDD NET61 NET72 VDD P18 W=1.64U L=0.18U
MP4 NET44 NETQ NET75 VDD P18 W=2.4U L=0.18U
MP5 VDD NET65 NET75 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET44 VDD P18 W=2.4U L=0.18U
MP0 NET78 NET24 NETQ VDD P18 W=0.6U L=0.18U
MP1 VDD NET61 NET81 VDD P18 W=3.36U L=0.18U
MN3 NET53 NETQ GND GND N18 W=1.18U L=0.18U
MN0 NETQ NET32 NET102 GND N18 W=0.3U L=0.18U
MN5 NET102 NET100 GND GND N18 W=0.3U L=0.18U
MN6 NETQ NET61 GND GND N18 W=0.72U L=0.18U
MN2 NET53 K GND GND N18 W=1.18U L=0.18U
MN4 NET68 NET33 GND GND N18 W=1.86U L=0.19U
MN1 NET75 NET65 NET53 GND N18 W=1.18U L=0.18U
XI18 NET65 NETQ J ND2G PW=0.51U NW=0.42U
XI9 NET68 NETQ NET24 NET32 TG1G NW=1.18U PW=1.18U
XI6 NET75 NET33 NET32 NET24 TG1G NW=0.6U PW=0.6U
.ENDS FFJKSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSHD2X                                                            *
* LAST TIME SAVED: MAR 13 14:19:05 2003                                       *
*******************************************************************************
.SUBCKT FFJKSHD2X Q QN CK J K SN
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI21 NET60 SN IVG PW=0.64U NW=0.42U
XI5 QN NET113 IVG PW=2.4U NW=1.6U
XI13 NET69 NET64 IVG PW=0.84U NW=0.42U
XI10 NET113 NETQ IVG PW=0.84U NW=0.56U
XI4 NET64 CK IVG PW=1.2U NW=0.6U
XI9 NET109 NETQ NET69 NET64 TG1G NW=1.1U PW=1.1U
XI6 NET35 NET71 NET64 NET69 TG1G NW=0.42U PW=0.42U
XI32 NET71 NET109 NET69 NET64 TRIIVG NW=0.3U PW=0.42U
MP1 VDD NET60 NET91 VDD P18 W=1.68U L=0.18U
MP4 NET36 NETQ NET35 VDD P18 W=1.66U L=0.18U
MP0 NET85 NET69 NETQ VDD P18 W=0.6U L=0.18U
MP7 NET88 NET113 NET85 VDD P18 W=0.6U L=0.18U
MP6 NET91 NET71 NET109 VDD P18 W=1.68U L=0.18U
MP5 VDD NET66 NET35 VDD P18 W=1.08U L=0.18U
MP2 VDD NET60 NET88 VDD P18 W=1.68U L=0.18U
MP3 VDD K NET36 VDD P18 W=1.66U L=0.18U
MN0 NETQ NET64 NET115 GND N18 W=0.3U L=0.18U
MN6 NETQ NET60 GND GND N18 W=0.72U L=0.18U
MN4 NET109 NET71 GND GND N18 W=0.9U L=0.18U
MN3 NET48 NETQ GND GND N18 W=0.9U L=0.18U
MN5 NET115 NET113 GND GND N18 W=0.3U L=0.18U
MN2 NET48 K GND GND N18 W=0.9U L=0.18U
MN1 NET35 NET66 NET48 GND N18 W=0.9U L=0.18U
XI18 NET66 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKSHD1X                                                            *
* LAST TIME SAVED: MAR 13 14:16:24 2003                                       *
*******************************************************************************
.SUBCKT FFJKSHD1X Q QN CK J K SN
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET138 CK IVG PW=0.84U NW=0.42U
XI21 NET56 SN IVG PW=0.64U NW=0.42U
XI13 NET67 NET138 IVG PW=0.6U NW=0.3U
XI5 QN NET105 IVG PW=1.2U NW=0.8U
XI10 NET105 NETQ IVG PW=0.64U NW=0.42U
XI6 NET42 NET69 NET138 NET67 TG1G NW=0.42U PW=0.42U
XI9 NET73 NETQ NET67 NET138 TG1G NW=0.7U PW=0.7U
XI31 NET69 NET73 NET67 NET138 TRIIVG NW=0.3U PW=0.42U
MP4 NET43 NETQ NET42 VDD P18 W=1.6U L=0.18U
MP5 VDD NET64 NET42 VDD P18 W=0.96U L=0.18U
MP1 VDD NET56 NET80 VDD P18 W=1.6U L=0.18U
MP3 VDD K NET43 VDD P18 W=1.6U L=0.18U
MP0 VDD NET56 NET83 VDD P18 W=1U L=0.18U
MP7 NET83 NET105 NET77 VDD P18 W=0.6U L=0.18U
MP6 NET80 NET69 NET73 VDD P18 W=1.6U L=0.18U
MP2 NET77 NET67 NETQ VDD P18 W=0.6U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.8U L=0.18U
MN6 NETQ NET56 GND GND N18 W=0.42U L=0.18U
MN0 NETQ NET138 NET107 GND N18 W=0.3U L=0.18U
MN5 NET107 NET105 GND GND N18 W=0.3U L=0.18U
MN4 NET73 NET69 GND GND N18 W=0.86U L=0.18U
MN2 NET52 K GND GND N18 W=0.8U L=0.18U
MN1 NET42 NET64 NET52 GND N18 W=0.8U L=0.18U
XI18 NET64 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKRHDLX                                                            *
* LAST TIME SAVED: NOV 25 17:36:57 2003                                       *
*******************************************************************************
.SUBCKT FFJKRHDLX Q QN CK J K RN
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET112 NETQ IVG PW=0.42U NW=0.3U
XI5 QN NET112 IVG PW=0.64U NW=0.42U
XI13 NET67 NET164 IVG PW=0.6U NW=0.3U
XI4 NET164 CK IVG PW=0.84U NW=0.42U
XI9 NET120 NETQ NET67 NET164 TG1G NW=0.7U PW=0.7U
XI6 NET39 NET69 NET164 NET67 TG1G NW=0.42U PW=0.42U
XI33 NET69 NET120 NET67 NET164 TRIIVG NW=0.3U PW=0.42U
MP0 NET99 NET67 NETQ VDD P18 W=0.45U L=0.18U
MP8 VDD RN NETQ VDD P18 W=0.64U L=0.18U
MP6 VDD NET112 NET99 VDD P18 W=0.45U L=0.18U
MP9 VDD NET69 NET120 VDD P18 W=0.88U L=0.18U
MP4 NET40 NETQ NET39 VDD P18 W=1.2U L=0.18U
MP5 VDD NET62 NET39 VDD P18 W=0.72U L=0.18U
MP3 VDD K NET40 VDD P18 W=1.2U L=0.18U
MN5 NET126 RN GND GND N18 W=0.6U L=0.18U
MN0 NET123 RN GND GND N18 W=0.77U L=0.18U
MN4 NET120 NET69 NET123 GND N18 W=0.77U L=0.18U
MN7 NETQ NET164 NET114 GND N18 W=0.3U L=0.18U
MN8 NET114 NET112 NET126 GND N18 W=0.3U L=0.18U
MN3 NET52 NETQ GND GND N18 W=0.6U L=0.18U
MN2 NET52 K GND GND N18 W=0.6U L=0.18U
MN1 NET39 NET62 NET52 GND N18 W=0.6U L=0.18U
XI18 NET62 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKRHD4X                                                            *
* LAST TIME SAVED: NOV 25 17:34:19 2003                                       *
*******************************************************************************
.SUBCKT FFJKRHD4X Q QN CK J K RN
XI12 Q NET214 IVG PW=4.8U NW=3.2U
XI10 NET242 NET214 IVG PW=1.68U NW=1.14U
XI5 QN NET242 IVG PW=4.8U NW=3.2U
XI13 NET189 NET190 IVG PW=0.96U NW=0.48U
XI4 NET190 CK IVG PW=1.2U NW=0.6U
XI9 NET247 NET214 NET189 NET190 TG1G NW=1.18U PW=1.18U
XI6 NET198 NET191 NET190 NET189 TG1G NW=0.6U PW=0.6U
XI33 NET191 NET247 NET189 NET190 TRIIVG NW=0.3U PW=0.42U
MP4 NET199 NET214 NET198 VDD P18 W=2.4U L=0.18U
MP5 VDD NET256 NET198 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET199 VDD P18 W=2.4U L=0.18U
MP0 NET217 NET189 NET214 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET214 VDD P18 W=1.1U L=0.18U
MP6 VDD NET191 NET247 VDD P18 W=2.52U L=0.18U
MP1 VDD NET242 NET217 VDD P18 W=0.45U L=0.18U
MN2 NET229 K GND GND N18 W=1.18U L=0.18U
MN1 NET198 NET256 NET229 GND N18 W=1.18U L=0.18U
MN3 NET229 NET214 GND GND N18 W=1.18U L=0.18U
MN7 NET238 RN GND GND N18 W=2.3U L=0.18U
MN8 NET244 NET242 NET253 GND N18 W=0.3U L=0.18U
MN0 NET247 NET191 NET238 GND N18 W=2.3U L=0.18U
MN4 NET214 NET190 NET244 GND N18 W=0.3U L=0.18U
MN5 NET253 RN GND GND N18 W=0.8U L=0.18U
XI18 NET256 NET214 J ND2G PW=0.51U NW=0.42U
.ENDS FFJKRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKRHD2X                                                            *
* LAST TIME SAVED: NOV 25 17:30:53 2003                                       *
*******************************************************************************
.SUBCKT FFJKRHD2X Q QN CK J K RN
XI12 Q NET257 IVG PW=2.4U NW=1.6U
XI10 NET116 NET257 IVG PW=0.84U NW=0.56U
XI5 QN NET116 IVG PW=2.4U NW=1.6U
XI36 NET65 NET63 IVG PW=0.84U NW=0.42U
XI4 NET63 CK IVG PW=1.2U NW=0.6U
XI9 NET121 NET257 NET65 NET63 TG1G NW=1.1U PW=1.1U
XI6 NET45 NET70 NET63 NET65 TG1G NW=0.42U PW=0.42U
XI33 NET70 NET121 NET65 NET63 TRIIVG NW=0.3U PW=0.42U
MP1 VDD NET116 NET97 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET257 VDD P18 W=0.64U L=0.18U
MP4 NET109 NET257 NET45 VDD P18 W=1.66U L=0.18U
MP5 VDD NET62 NET45 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET109 VDD P18 W=1.66U L=0.18U
MP6 VDD NET70 NET121 VDD P18 W=1.28U L=0.18U
MP0 NET97 NET65 NET257 VDD P18 W=0.45U L=0.18U
MN3 NET55 NET257 GND GND N18 W=0.9U L=0.18U
MN4 NET121 NET70 NET124 GND N18 W=1.12U L=0.18U
MN5 NET118 NET116 NET115 GND N18 W=0.3U L=0.18U
MN7 NET115 RN GND GND N18 W=0.6U L=0.18U
MN8 NET257 NET63 NET118 GND N18 W=0.3U L=0.18U
MN0 NET124 RN GND GND N18 W=1.12U L=0.18U
MN2 NET55 K GND GND N18 W=0.9U L=0.18U
MN1 NET45 NET62 NET55 GND N18 W=0.9U L=0.18U
XI18 NET62 NET257 J ND2G PW=0.51U NW=0.42U
.ENDS FFJKRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKRHD1X                                                            *
* LAST TIME SAVED: NOV 13 10:47:44 2003                                       *
*******************************************************************************
.SUBCKT FFJKRHD1X Q QN CK J K RN
XI9 NET135 NETQ NET59 NET74 TG1G NW=0.7U PW=0.7U
XI6 NET45 NET61 NET74 NET59 TG1G NW=0.42U PW=0.42U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NET115 NETQ IVG PW=0.64U NW=0.42U
XI13 NET59 NET74 IVG PW=0.6U NW=0.3U
XI4 NET74 CK IVG PW=0.84U NW=0.42U
XI5 QN NET115 IVG PW=1.2U NW=0.8U
XI34 NET61 NET135 NET59 NET74 TRIIVG NW=0.3U PW=0.42U
MP4 NET107 NETQ NET45 VDD P18 W=1.6U L=0.18U
MP5 VDD NET58 NET45 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET107 VDD P18 W=1.6U L=0.18U
MP0 VDD NET115 NET87 VDD P18 W=0.45U L=0.18U
MP2 NET87 NET59 NETQ VDD P18 W=0.45U L=0.18U
MP8 VDD RN NETQ VDD P18 W=0.64U L=0.18U
MP9 VDD NET61 NET135 VDD P18 W=1.28U L=0.18U
MN3 NET55 NETQ GND GND N18 W=0.8U L=0.18U
MN0 NETQ NET74 NET117 GND N18 W=0.3U L=0.18U
MN2 NET55 K GND GND N18 W=0.8U L=0.18U
MN7 NET129 RN GND GND N18 W=1.06U L=0.18U
MN4 NET117 NET115 NET114 GND N18 W=0.3U L=0.18U
MN1 NET45 NET58 NET55 GND N18 W=0.8U L=0.18U
MN5 NET114 RN GND GND N18 W=0.6U L=0.18U
MN8 NET135 NET61 NET129 GND N18 W=1.06U L=0.18U
XI33 NET58 NETQ J ND2G PW=0.51U NW=0.42U
.ENDS FFJKRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKHDLX                                                             *
* LAST TIME SAVED: MAR  4 15:37:37 2003                                       *
*******************************************************************************
.SUBCKT FFJKHDLX Q QN CK J K
MP4 NET34 NETQ NET100 VDD P18 W=1.2U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=0.72U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.2U L=0.18U
MN2 NET101 K GND GND N18 W=0.6U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.6U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.6U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.52U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI6 NET100 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET32 NET96 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=0.64U NW=0.42U
XI4 NET96 CK IVG PW=0.84U NW=0.42U
.ENDS FFJKHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKHD4X                                                             *
* LAST TIME SAVED: MAR  4 15:37:21 2003                                       *
*******************************************************************************
.SUBCKT FFJKHD4X Q QN CK J K
MP4 NET34 NETQ NET100 VDD P18 W=2.4U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=1.42U L=0.18U
MP3 VDD K NET34 VDD P18 W=2.4U L=0.18U
MN2 NET101 K GND GND N18 W=1.18U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=1.18U L=0.18U
MN3 NET101 NETQ GND GND N18 W=1.18U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI6 NET100 NET33 NET96 NET32 TG1G NW=0.6U PW=0.6U
XI9 NET46 NETQ NET32 NET96 TG1G NW=1.18U PW=1.18U
XI7 NET46 NET33 IVG PW=3.44U NW=2.44U
XI13 NET32 NET96 IVG PW=0.96U NW=0.48U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.68U NW=1.14U
XI5 QN NETQN IVG PW=4.8U NW=3.2U
XI4 NET96 CK IVG PW=1.2U NW=0.6U
.ENDS FFJKHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKHD2X                                                             *
* LAST TIME SAVED: MAR  4 15:37:03 2003                                       *
*******************************************************************************
.SUBCKT FFJKHD2X Q QN CK J K
MP4 NET34 NETQ NET100 VDD P18 W=1.66U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=1.08U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.66U L=0.18U
MN2 NET101 K GND GND N18 W=0.9U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.9U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.9U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI6 NET100 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=1.1U PW=1.1U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI13 NET32 NET96 IVG PW=0.84U NW=0.42U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 QN NETQN IVG PW=2.4U NW=1.6U
XI4 NET96 CK IVG PW=1.2U NW=0.6U
.ENDS FFJKHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFJKHD1X                                                             *
* LAST TIME SAVED: DEC  1 15:38:21 2003                                       *
*******************************************************************************
.SUBCKT FFJKHD1X Q QN CK J K
MP4 NET34 NETQ NET100 VDD P18 W=1.6U L=0.18U
MP5 VDD NET52 NET100 VDD P18 W=0.96U L=0.18U
MP3 VDD K NET34 VDD P18 W=1.6U L=0.18U
MN2 NET101 K GND GND N18 W=0.8U L=0.18U
MN1 NET100 NET52 NET101 GND N18 W=0.8U L=0.18U
MN3 NET101 NETQ GND GND N18 W=0.8U L=0.18U
XI18 NET52 NETQ J ND2G PW=0.51U NW=0.42U
XI17 NET33 NET46 NET32 NET96 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET96 NET32 TRIIVG NW=0.3U PW=0.42U
XI6 NET100 NET33 NET96 NET32 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET32 NET96 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET32 NET96 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 QN NETQN IVG PW=1.2U NW=0.8U
XI4 NET96 CK IVG PW=0.84U NW=0.42U
.ENDS FFJKHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDQHDLX                                                            *
* LAST TIME SAVED: DEC  1 14:53:18 2003                                       *
*******************************************************************************
.SUBCKT FFEDQHDLX Q CK D E
XI21 NET42 NETQN NET61 E TRIIVG NW=0.32U PW=0.48U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET33 NET42 NET32 NET24 TRIIVG NW=0.45U PW=0.51U
XI22 NET42 D E NET61 TRIIVG NW=0.32U PW=0.48U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFEDQHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDQHD4X                                                            *
* LAST TIME SAVED: DEC  1 14:52:43 2003                                       *
*******************************************************************************
.SUBCKT FFEDQHD4X Q CK D E
XI21 NET42 NETQN NET61 E TRIIVG NW=0.6U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET33 NET42 NET32 NET24 TRIIVG NW=1U PW=1.17U
XI22 NET42 D E NET61 TRIIVG NW=0.6U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.81U NW=1.81U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
.ENDS FFEDQHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDQHD2X                                                            *
* LAST TIME SAVED: DEC  1 14:52:14 2003                                       *
*******************************************************************************
.SUBCKT FFEDQHD2X Q CK D E
XI21 NET42 NETQN NET61 E TRIIVG NW=0.42U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET33 NET42 NET32 NET24 TRIIVG NW=0.51U PW=0.69U
XI22 NET42 D E NET61 TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFEDQHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDQHD1X                                                            *
* LAST TIME SAVED: DEC  1 14:51:44 2003                                       *
*******************************************************************************
.SUBCKT FFEDQHD1X Q CK D E
XI21 NET42 NETQN NET61 E TRIIVG NW=0.42U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI23 NET33 NET42 NET32 NET24 TRIIVG NW=0.42U PW=0.64U
XI22 NET42 D E NET61 TRIIVG NW=0.42U PW=0.64U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFEDQHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDHDLX                                                             *
* LAST TIME SAVED: DEC  1 14:55:23 2003                                       *
*******************************************************************************
.SUBCKT FFEDHDLX Q QN CK D E
XI21 NET42 NETQ NET61 E TRIIVG NW=0.54U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET42 D E NET61 TRIIVG NW=0.54U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET42 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFEDHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDHD4X                                                             *
* LAST TIME SAVED: DEC  1 14:54:59 2003                                       *
*******************************************************************************
.SUBCKT FFEDHD4X Q QN CK D E
XI21 NET42 NETQ NET61 E TRIIVG NW=0.9U PW=1.5U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET42 D E NET61 TRIIVG NW=0.9U PW=1.5U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET42 NET33 NET32 NET24 TG1G NW=0.7U PW=0.7U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=2.52U NW=1.68U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
.ENDS FFEDHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDHD2X                                                             *
* LAST TIME SAVED: DEC  1 14:54:12 2003                                       *
*******************************************************************************
.SUBCKT FFEDHD2X Q QN CK D E
XI21 NET42 NETQ NET61 E TRIIVG NW=0.54U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET42 D E NET61 TRIIVG NW=0.54U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET42 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFEDHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDHD1X                                                             *
* LAST TIME SAVED: DEC  1 14:53:44 2003                                       *
*******************************************************************************
.SUBCKT FFEDHD1X Q QN CK D E
XI21 NET42 NETQ NET61 E TRIIVG NW=0.54U PW=0.9U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI22 NET42 D E NET61 TRIIVG NW=0.54U PW=0.9U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET42 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI20 NET61 E IVG PW=0.42U NW=0.3U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFEDHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDCRHDLX                                                           *
* LAST TIME SAVED: MAR  4 15:07:48 2003                                       *
*******************************************************************************
.SUBCKT FFEDCRHDLX Q QN CK D E RN
XI18 NET63 RN NET54 ND2G PW=0.6U NW=0.5U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI20 NETQN NET54 NET65 E TG1G NW=0.42U PW=0.42U
XI19 D NET54 E NET65 TG1G NW=0.42U PW=0.42U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=0.64U NW=0.42U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFEDCRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDCRHD4X                                                           *
* LAST TIME SAVED: MAR  4 15:07:27 2003                                       *
*******************************************************************************
.SUBCKT FFEDCRHD4X Q QN CK D E RN
XI18 NET63 RN NET54 ND2G PW=1.47U NW=1.18U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI20 NETQN NET54 NET65 E TG1G NW=0.7U PW=0.7U
XI19 D NET54 E NET65 TG1G NW=0.7U PW=0.7U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.6U PW=0.6U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.18U PW=1.18U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=3.44U NW=2.3U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI12 QN NETQN IVG PW=4.8U NW=3.2U
XI10 NETQ NETQN IVG PW=1.68U NW=1.14U
XI5 Q NETQ IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFEDCRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDCRHD2X                                                           *
* LAST TIME SAVED: MAR  4 15:07:10 2003                                       *
*******************************************************************************
.SUBCKT FFEDCRHD2X Q QN CK D E RN
XI18 NET63 RN NET54 ND2G PW=0.96U NW=0.8U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI20 NETQN NET54 NET65 E TG1G NW=0.6U PW=0.6U
XI19 D NET54 E NET65 TG1G NW=0.6U PW=0.6U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFEDCRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFEDCRHD1X                                                           *
* LAST TIME SAVED: MAR  4 15:06:51 2003                                       *
*******************************************************************************
.SUBCKT FFEDCRHD1X Q QN CK D E RN
XI18 NET63 RN NET54 ND2G PW=0.66U NW=0.55U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI20 NETQN NET54 NET65 E TG1G NW=0.6U PW=0.6U
XI19 D NET54 E NET65 TG1G NW=0.6U PW=0.6U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI21 NET65 E IVG PW=0.64U NW=0.42U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=1.2U NW=0.8U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFEDCRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSRHDLX                                                            *
* LAST TIME SAVED: DEC  1 15:02:30 2003                                       *
*******************************************************************************
.SUBCKT FFDSRHDLX Q QN CK D RN SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.38U PW=0.64U
XI21 NET53 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 QN NET95 IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.64U NW=0.42U
XI5 Q NET60 IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN0 NET79 NET53 GND GND N18 W=0.54U L=0.18U
MN6 NET95 SN NET79 GND N18 W=0.54U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=0.72U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=0.72U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=1.1U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET122 NET65 VDD P18 W=1.1U L=0.18U
XI9 NET65 NET95 NET24 NET32 TG1G NW=0.5U PW=0.5U
.ENDS FFDSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSRHD4X                                                            *
* LAST TIME SAVED: DEC 27 23:13:56 2003                                       *
*******************************************************************************
.SUBCKT FFDSRHD4X Q QN CK D RN SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.78U PW=1.32U
XI21 NET53 RN IVG PW=1.5U NW=1U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NET95 IVG PW=4.8U NW=3.2U
XI10 NET60 NET95 IVG PW=1.77U NW=1.18U
XI5 Q NET60 IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN0 NET79 NET53 GND GND N18 W=0.92U L=0.18U
MN6 NET95 SN NET79 GND N18 W=0.92U L=0.18U
MN5 NET59 SN GND GND N18 W=0.8U L=0.18U
MN3 NET68 SN GND GND N18 W=2.16U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=2.16U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=3.3U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1.68U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET95 VDD P18 W=1.1U L=0.18U
MP6 NET89 NET122 NET65 VDD P18 W=3.3U L=0.18U
XI9 NET65 NET95 NET24 NET32 TG1G NL=0.19U NW=1.35U PL=0.19U PW=1.35U
.ENDS FFDSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSRHD2X                                                            *
* LAST TIME SAVED: DEC  1 15:01:58 2003                                       *
*******************************************************************************
.SUBCKT FFDSRHD2X Q QN CK D RN SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.54U PW=0.96U
XI21 NET53 RN IVG PW=0.81U NW=0.54U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NET95 IVG PW=2.4U NW=1.6U
XI10 NET60 NET95 IVG PW=0.84U NW=0.56U
XI5 Q NET60 IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN0 NET79 NET53 GND GND N18 W=0.54U L=0.18U
MN6 NET95 SN NET79 GND N18 W=0.54U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.57U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=1.57U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=2.25U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=0.86U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET122 NET65 VDD P18 W=2.25U L=0.18U
XI9 NET65 NET95 NET24 NET32 TG1G NW=1.1U PW=1.1U
.ENDS FFDSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSRHD1X                                                            *
* LAST TIME SAVED: DEC  1 15:01:43 2003                                       *
*******************************************************************************
.SUBCKT FFDSRHD1X Q QN CK D RN SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.42U PW=0.84U
XI21 NET53 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NET95 IVG PW=1.2U NW=0.8U
XI10 NET60 NET95 IVG PW=0.64U NW=0.42U
XI5 Q NET60 IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN0 NET79 NET53 GND GND N18 W=0.54U L=0.18U
MN6 NET95 SN NET79 GND N18 W=0.54U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.1U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=1.1U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=1.68U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET122 NET65 VDD P18 W=1.68U L=0.18U
XI9 NET65 NET95 NET24 NET32 TG1G NW=0.7U PW=0.7U
.ENDS FFDSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSHDLX                                                             *
* LAST TIME SAVED: DEC  1 15:03:32 2003                                       *
*******************************************************************************
.SUBCKT FFDSHDLX Q QN CK D SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.38U PW=0.64U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 QN NET105 IVG PW=0.64U NW=0.42U
XI10 NET60 NET105 IVG PW=0.64U NW=0.42U
XI5 Q NET60 IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET105 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=0.72U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=0.72U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET105 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET105 VDD P18 W=0.64U L=0.18U
MP6 VDD NET122 NET65 VDD P18 W=0.84U L=0.18U
XI9 NET65 NET105 NET24 NET32 TG1G NW=0.5U PW=0.5U
.ENDS FFDSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSHD4X                                                             *
* LAST TIME SAVED: DEC  1 15:03:17 2003                                       *
*******************************************************************************
.SUBCKT FFDSHD4X Q QN CK D SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.78U PW=1.32U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NET105 IVG PW=4.8U NW=3.2U
XI10 NET60 NET105 IVG PW=1.77U NW=1.18U
XI5 Q NET60 IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
MN1 NET105 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 SN GND GND N18 W=0.8U L=0.18U
MN3 NET68 SN GND GND N18 W=2.16U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=2.16U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET105 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET105 VDD P18 W=1.1U L=0.18U
MP6 VDD NET122 NET65 VDD P18 W=2.52U L=0.18U
XI9 NET65 NET105 NET24 NET32 TG1G NW=1.35U PW=1.35U
.ENDS FFDSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSHD2X                                                             *
* LAST TIME SAVED: DEC 27 23:06:28 2003                                       *
*******************************************************************************
.SUBCKT FFDSHD2X Q QN CK D SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.54U PW=0.96U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NET105 IVG PW=2.4U NW=1.6U
XI10 NET60 NET105 IVG PW=0.84U NW=0.56U
XI5 Q NET60 IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
MN1 NET105 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.57U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=1.57U L=0.19U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET105 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET105 VDD P18 W=0.91U L=0.18U
MP6 VDD NET122 NET65 VDD P18 W=1.72U L=0.18U
XI9 NET65 NET105 NET24 NET32 TG1G NW=1.1U PW=1.1U
.ENDS FFDSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDSHD1X                                                             *
* LAST TIME SAVED: DEC  1 15:02:46 2003                                       *
*******************************************************************************
.SUBCKT FFDSHD1X Q QN CK D SN
XI32 NET122 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET122 D NET32 NET24 TRIIVG NW=0.42U PW=0.84U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NET105 IVG PW=1.2U NW=0.8U
XI10 NET60 NET105 IVG PW=0.64U NW=0.42U
XI5 Q NET60 IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET105 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.06U L=0.18U
MN2 NET65 NET122 NET68 GND N18 W=1.06U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET105 VDD P18 W=0.45U L=0.18U
MP8 VDD SN NET105 VDD P18 W=0.64U L=0.18U
MP6 VDD NET122 NET65 VDD P18 W=1.28U L=0.18U
XI9 NET65 NET105 NET24 NET32 TG1G NW=0.7U PW=0.7U
.ENDS FFDSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDRHDLX                                                             *
* LAST TIME SAVED: DEC  1 15:04:48 2003                                       *
*******************************************************************************
.SUBCKT FFDRHDLX Q QN CK D RN
MN1 NET70 NET32 NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 NET36 GND GND N18 W=0.3U L=0.18U
MN3 NET62 NET33 GND GND N18 W=0.56U L=0.18U
MN6 NET70 NET79 GND GND N18 W=0.42U L=0.18U
MP1 VDD NET79 NET56 VDD P18 W=1.1U L=0.18U
MP5 VDD NET79 NET53 VDD P18 W=1U L=0.18U
MP7 NET53 NET36 NET59 VDD P18 W=0.42U L=0.18U
MP6 NET56 NET33 NET62 VDD P18 W=1.1U L=0.18U
MP4 NET59 NET24 NET70 VDD P18 W=0.42U L=0.18U
XI29 NET33 NET62 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET32 NET24 TRIIVG NW=0.38U PW=0.64U
XI9 NET62 NET70 NET24 NET32 TG1G NW=0.5U PW=0.5U
XI12 QN NET70 IVG PW=0.64U NW=0.42U
XI10 NET36 NET70 IVG PW=0.64U NW=0.42U
XI5 Q NET36 IVG PW=0.64U NW=0.42U
XI21 NET79 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDRHD4X                                                             *
* LAST TIME SAVED: DEC  1 15:04:31 2003                                       *
*******************************************************************************
.SUBCKT FFDRHD4X Q QN CK D RN
MN1 NET70 NET32 NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 NET36 GND GND N18 W=0.3U L=0.18U
MN3 NET62 NET33 GND GND N18 W=1.68U L=0.18U
MN6 NET70 NET79 GND GND N18 W=0.72U L=0.18U
MP1 VDD NET79 NET56 VDD P18 W=3.3U L=0.18U
MP5 VDD NET79 NET53 VDD P18 W=1.68U L=0.18U
MP7 NET53 NET36 NET59 VDD P18 W=0.42U L=0.18U
MP6 NET56 NET33 NET62 VDD P18 W=3.3U L=0.18U
MP4 NET59 NET24 NET70 VDD P18 W=0.42U L=0.18U
XI29 NET33 NET62 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET32 NET24 TRIIVG NW=0.78U PW=1.32U
XI9 NET62 NET70 NET24 NET32 TG1G NW=1.36U PW=1.36U
XI12 QN NET70 IVG PW=4.8U NW=3.2U
XI10 NET36 NET70 IVG PW=1.77U NW=1.18U
XI5 Q NET36 IVG PW=4.8U NW=3.2U
XI21 NET79 RN IVG PW=1.5U NW=1U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
.ENDS FFDRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDRHD2X                                                             *
* LAST TIME SAVED: DEC  1 15:04:16 2003                                       *
*******************************************************************************
.SUBCKT FFDRHD2X Q QN CK D RN
MN1 NET70 NET32 NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 NET36 GND GND N18 W=0.3U L=0.18U
MN3 NET62 NET33 GND GND N18 W=1.22U L=0.18U
MN6 NET70 NET79 GND GND N18 W=0.42U L=0.18U
MP1 VDD NET79 NET56 VDD P18 W=2.25U L=0.18U
MP5 VDD NET79 NET53 VDD P18 W=0.86U L=0.18U
MP7 NET53 NET36 NET59 VDD P18 W=0.42U L=0.18U
MP6 NET56 NET33 NET62 VDD P18 W=2.25U L=0.18U
MP4 NET59 NET24 NET70 VDD P18 W=0.42U L=0.18U
XI29 NET33 NET62 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET32 NET24 TRIIVG NW=0.54U PW=0.96U
XI9 NET62 NET70 NET24 NET32 TG1G NW=1.1U PW=1.1U
XI12 QN NET70 IVG PW=2.4U NW=1.6U
XI10 NET36 NET70 IVG PW=0.84U NW=0.56U
XI5 Q NET36 IVG PW=2.4U NW=1.6U
XI21 NET79 RN IVG PW=0.81U NW=0.54U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFDRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDRHD1X                                                             *
* LAST TIME SAVED: DEC  1 15:03:51 2003                                       *
*******************************************************************************
.SUBCKT FFDRHD1X Q QN CK D RN
MN1 NET70 NET32 NET38 GND N18 W=0.3U L=0.18U
MN5 NET38 NET36 GND GND N18 W=0.3U L=0.18U
MN3 NET62 NET33 GND GND N18 W=0.86U L=0.18U
MN6 NET70 NET79 GND GND N18 W=0.42U L=0.18U
MP1 VDD NET79 NET56 VDD P18 W=1.68U L=0.18U
MP5 VDD NET79 NET53 VDD P18 W=1U L=0.18U
MP7 NET53 NET36 NET59 VDD P18 W=0.42U L=0.18U
MP6 NET56 NET33 NET62 VDD P18 W=1.68U L=0.18U
MP4 NET59 NET24 NET70 VDD P18 W=0.42U L=0.18U
XI29 NET33 NET62 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET32 NET24 TRIIVG NW=0.42U PW=0.84U
XI9 NET62 NET70 NET24 NET32 TG1G NW=0.7U PW=0.7U
XI12 QN NET70 IVG PW=1.2U NW=0.8U
XI10 NET36 NET70 IVG PW=0.64U NW=0.42U
XI5 Q NET36 IVG PW=1.2U NW=0.8U
XI21 NET79 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSRHDLX                                                           *
* LAST TIME SAVED: DEC 13 14:31:00 2003                                       *
*******************************************************************************
.SUBCKT FFDQSRHDLX Q CK D RN SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.64U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=0.42U PW=0.64U
XI35 NET73 RN IVG PW=0.64U NW=0.42U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NET95 IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN0 NET65 SN NET86 GND N18 W=0.51U L=0.18U
MN7 NET86 NET73 GND GND N18 W=0.51U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=0.51U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=0.51U L=0.18U
MP0 VDD SN NET65 VDD P18 W=0.91U L=0.18U
MP1 VDD NET73 NET89 VDD P18 W=1.2U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP3 NET74 NET53 NET95 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET74 VDD P18 W=0.84U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=1.2U L=0.18U
.ENDS FFDQSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSRHD4X                                                           *
* LAST TIME SAVED: DEC 27 23:10:42 2003                                       *
*******************************************************************************
.SUBCKT FFDQSRHD4X Q CK D RN SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.65U PW=1.05U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=1.24U PW=1.86U
XI35 NET144 RN IVG PW=0.64U NW=0.42U
XI21 NET53 SN IVG PW=1.5U NW=1U PL=0.19U NL=0.18U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NET95 IVG PW=4.8U NW=3.2U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
MN0 NET65 SN NET90 GND N18 W=1.73U L=0.18U
MN7 NET90 NET144 GND GND N18 W=1.73U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.72U L=0.18U
MN5 NET59 RN GND GND N18 W=0.8U L=0.18U
MN3 NET68 SN GND GND N18 W=1.73U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.73U L=0.18U
MP1 VDD NET144 NET89 VDD P18 W=3.34U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1.68U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET65 VDD P18 W=2.55U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP3 NET74 NET53 NET95 VDD P18 W=1.44U L=0.19U
MP8 VDD RN NET74 VDD P18 W=1.44U L=0.19U
MP6 NET89 NET33 NET65 VDD P18 W=3.34U L=0.18U
.ENDS FFDQSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSRHD2X                                                           *
* LAST TIME SAVED: DEC 13 14:26:35 2003                                       *
*******************************************************************************
.SUBCKT FFDQSRHD2X Q CK D RN SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.45U PW=0.8U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=0.8U PW=1.2U
XI35 NET145 RN IVG PW=0.64U NW=0.42U
XI21 NET53 SN IVG PW=0.81U NW=0.54U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NET95 IVG PW=2.4U NW=1.6U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
MN0 NET65 SN NET87 GND N18 W=1.51U L=0.18U
MN7 NET87 NET145 GND GND N18 W=1.51U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.51U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.51U L=0.18U
MP0 VDD SN NET65 VDD P18 W=1.77U L=0.18U
MP1 VDD NET145 NET89 VDD P18 W=2.3U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=0.86U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP3 NET74 NET53 NET95 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET74 VDD P18 W=0.84U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=2.3U L=0.18U
.ENDS FFDQSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSRHD1X                                                           *
* LAST TIME SAVED: DEC 13 14:15:53 2003                                       *
*******************************************************************************
.SUBCKT FFDQSRHD1X Q CK D RN SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.75U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=0.56U PW=0.84U
XI35 NET73 RN IVG PW=0.64U NW=0.42U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET95 IVG PW=1.2U NW=0.8U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN0 NET65 SN NET86 GND N18 W=1.06U L=0.18U
MN7 NET86 NET73 GND GND N18 W=1.06U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN3 NET68 SN GND GND N18 W=1.06U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.06U L=0.18U
MP0 VDD SN NET65 VDD P18 W=1.28U L=0.18U
MP1 VDD NET73 NET89 VDD P18 W=1.6U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP3 NET74 NET53 NET95 VDD P18 W=0.84U L=0.18U
MP8 VDD RN NET74 VDD P18 W=0.84U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=1.6U L=0.18U
.ENDS FFDQSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSHDLX                                                            *
* LAST TIME SAVED: NOV 30 14:16:57 2003                                       *
*******************************************************************************
.SUBCKT FFDQSHDLX Q CK D SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.64U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=0.42U PW=0.64U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NET95 IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 GND GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN3 NET68 SN GND GND N18 W=0.51U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=0.51U L=0.18U
MP0 VDD SN NET65 VDD P18 W=0.45U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP6 VDD NET33 NET65 VDD P18 W=0.45U L=0.18U
.ENDS FFDQSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSHD4X                                                            *
* LAST TIME SAVED: DEC 27 18:40:00 2003                                       *
*******************************************************************************
.SUBCKT FFDQSHD4X Q CK D SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.65U PW=1.05U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=1.24U PW=1.86U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NET95 IVG PW=4.8U NW=3.2U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 GND GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.72U L=0.18U
MN3 NET68 SN GND GND N18 W=1.73U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.73U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1.68U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET65 VDD P18 W=2.55U L=0.19U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP6 VDD NET33 NET65 VDD P18 W=2.55U L=0.18U
.ENDS FFDQSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSHD2X                                                            *
* LAST TIME SAVED: DEC 27 18:40:38 2003                                       *
*******************************************************************************
.SUBCKT FFDQSHD2X Q CK D SN
XI32 NET33 NET65 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.45U PW=0.8U
XI34 NET95 NET65 NET24 NET32 TRIIVG NW=0.8U PW=1.2U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NET95 IVG PW=2.4U NW=1.6U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 GND GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN3 NET68 SN GND GND N18 W=1.51U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.51U L=0.18U
MP0 VDD SN NET65 VDD P18 W=1.77U L=0.19U
MP7 VDD NET53 NET77 VDD P18 W=0.86U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP6 VDD NET33 NET65 VDD P18 W=1.77U L=0.18U
.ENDS FFDQSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQSHD1X                                                            *
* LAST TIME SAVED: NOV 30 13:27:24 2003                                       *
*******************************************************************************
.SUBCKT FFDQSHD1X Q CK D SN
XI32 NET33 NET111 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.75U
XI34 NET95 NET111 NET24 NET32 TRIIVG NW=0.56U PW=0.84U
XI21 NET53 SN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET95 IVG PW=1.2U NW=0.8U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 GND GND N18 W=0.3U L=0.18U
MN6 NET95 NET53 GND GND N18 W=0.42U L=0.18U
MN8 NET68 SN GND GND N18 W=1.06U L=0.18U
MN2 NET111 NET33 NET68 GND N18 W=1.06U L=0.18U
MP0 VDD SN NET111 VDD P18 W=1.28U L=0.18U
MP7 VDD NET53 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP6 VDD NET33 NET111 VDD P18 W=1.28U L=0.18U
.ENDS FFDQSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQRHDLX                                                            *
* LAST TIME SAVED: NOV 30 14:08:14 2003                                       *
*******************************************************************************
.SUBCKT FFDQRHDLX Q CK D RN
XI32 NET33 NET87 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.64U
XI34 NET95 NET87 NET24 NET32 TRIIVG NW=0.42U PW=0.64U
XI35 NET53 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NET95 IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN7 NET87 NET53 GND GND N18 W=0.4U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN2 NET87 NET33 GND GND N18 W=0.4U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=0.6U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET33 NET87 VDD P18 W=0.6U L=0.18U
.ENDS FFDQRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQRHD4X                                                            *
* LAST TIME SAVED: NOV 30 14:04:57 2003                                       *
*******************************************************************************
.SUBCKT FFDQRHD4X Q CK D RN
XI32 NET33 NET90 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.65U PW=1.05U
XI34 NET95 NET90 NET24 NET32 TRIIVG NW=1.24U PW=1.86U
XI35 NET53 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NET95 IVG PW=4.8U NW=3.2U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
MN7 NET90 NET53 GND GND N18 W=1.35U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 RN GND GND N18 W=0.8U L=0.18U
MN2 NET90 NET33 GND GND N18 W=1.35U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=3.34U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET95 VDD P18 W=1.1U L=0.18U
MP6 NET89 NET33 NET90 VDD P18 W=3.34U L=0.18U
.ENDS FFDQRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQRHD2X                                                            *
* LAST TIME SAVED: NOV 30 14:02:03 2003                                       *
*******************************************************************************
.SUBCKT FFDQRHD2X Q CK D RN
XI32 NET33 NET87 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.45U PW=0.8U
XI34 NET95 NET87 NET24 NET32 TRIIVG NW=0.8U PW=1.2U
XI35 NET53 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NET95 IVG PW=2.4U NW=1.6U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
MN7 NET87 NET53 GND GND N18 W=1.18U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN2 NET87 NET33 GND GND N18 W=1.18U L=0.18U
MP1 VDD NET53 NET89 VDD P18 W=2.3U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET33 NET87 VDD P18 W=2.3U L=0.18U
.ENDS FFDQRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQRHD1X                                                            *
* LAST TIME SAVED: NOV 30 13:36:45 2003                                       *
*******************************************************************************
.SUBCKT FFDQRHD1X Q CK D RN
XI32 NET33 NET86 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.75U
XI34 NET95 NET86 NET24 NET32 TRIIVG NW=0.56U PW=0.84U
XI35 NET73 RN IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NET95 IVG PW=1.2U NW=0.8U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
MN7 NET86 NET73 GND GND N18 W=1.06U L=0.18U
MN1 NET95 NET32 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN5 NET59 RN GND GND N18 W=0.6U L=0.18U
MN2 NET86 NET33 GND GND N18 W=1.06U L=0.18U
MP1 VDD NET73 NET89 VDD P18 W=1.6U L=0.18U
MP5 VDD NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET24 NET95 VDD P18 W=0.45U L=0.18U
MP8 VDD RN NET95 VDD P18 W=0.84U L=0.18U
MP6 NET89 NET33 NET86 VDD P18 W=1.6U L=0.18U
.ENDS FFDQRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQHDLX                                                             *
* LAST TIME SAVED: NOV 24 16:10:34 2003                                       *
*******************************************************************************
.SUBCKT FFDQHDLX Q CK D
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.64U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET43 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI18 NET43 NET46 IVG PW=0.91U NW=0.4U
XI7 NET46 NET33 IVG PW=0.46U NW=0.41U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI12 Q NETQ IVG PW=0.64U NW=0.42U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDQHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQHD4X                                                             *
* LAST TIME SAVED: NOV 24 15:29:50 2003                                       *
*******************************************************************************
.SUBCKT FFDQHD4X Q CK D
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI19 NET33 D NET32 NET24 TRIIVG NW=0.65U PW=1.05U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET45 NETQ NET24 NET32 TG1G NW=1.2U PW=1.2U
XI7 NET46 NET33 IVG PW=1.05U NW=0.96U
XI18 NET45 NET46 IVG PW=2.55U NW=1.35U PL=0.18U NL=0.19U
XI13 NET24 NET32 IVG PW=0.9U NW=0.3U
XI12 Q NETQ IVG PW=4.8U NW=3.2U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.75U
.ENDS FFDQHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQHD2X                                                             *
* LAST TIME SAVED: NOV 24 13:16:58 2003                                       *
*******************************************************************************
.SUBCKT FFDQHD2X Q CK D
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET32 NET24 TRIIVG NW=0.45U PW=0.8U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 NET75 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI19 NET75 NET46 IVG PW=1.76U NW=1.18U
XI7 NET46 NET33 IVG PW=0.81U NW=0.72U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 Q NETQ IVG PW=2.4U NW=1.6U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFDQHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDQHD1X                                                             *
* LAST TIME SAVED: DEC  1 15:05:25 2003                                       *
*******************************************************************************
.SUBCKT FFDQHD1X Q CK D
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET32 NET24 TRIIVG NW=0.3U PW=0.75U
XI11 NETQ NET9 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET45 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI19 NET45 NET46 IVG PW=1.28U NW=0.86U
XI7 NET46 NET33 IVG PW=0.58U NW=0.48U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 Q NETQ IVG PW=1.2U NW=0.8U
XI10 NET9 NETQ IVG PW=0.42U NW=0.3U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDQHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSRHDLX                                                           *
* LAST TIME SAVED: DEC  1 15:07:39 2003                                       *
*******************************************************************************
.SUBCKT FFDNSRHDLX Q QN CKN D RN SN
XI32 NET33 NET65 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NET95 IVG PW=0.64U NW=0.42U
XI34 NET128 RN IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.42U NW=0.3U
XI5 Q NET60 IVG PW=0.64U NW=0.42U
XI4 NET32 CKN IVG PW=0.9U NW=0.3U
MN1 NET95 NET24 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 SN NET83 GND N18 W=0.58U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN0 NET83 NET128 GND GND N18 W=0.58U L=0.18U
MN3 NET68 SN GND GND N18 W=0.64U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=0.64U L=0.18U
MP1 VDD NET128 NET89 VDD P18 W=1.1U L=0.18U
MP7 VDD NET128 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET32 NET95 VDD P18 W=0.45U L=0.18U
MP3 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=1.1U L=0.18U
XI9 NET65 NET95 NET32 NET24 TG1G NW=0.5U PW=0.5U
.ENDS FFDNSRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSRHD4X                                                           *
* LAST TIME SAVED: DEC 27 23:12:38 2003                                       *
*******************************************************************************
.SUBCKT FFDNSRHD4X Q QN CKN D RN SN
XI32 NET33 NET65 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET24 NET32 TRIIVG NW=0.45U PW=1.62U
XI13 NET24 NET32 IVG PW=0.3U NW=0.48U
XI12 QN NET95 IVG PW=4.8U NW=3.2U
XI34 NET128 RN IVG PW=1.5U NW=1U
XI10 NET60 NET95 IVG PW=1.77U NW=1.18U
XI5 Q NET60 IVG PW=4.8U NW=3.2U
XI4 NET32 CKN IVG PW=1.44U NW=0.3U
MN1 NET95 NET24 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 SN NET83 GND N18 W=0.92U L=0.18U
MN5 NET59 SN GND GND N18 W=0.8U L=0.18U
MN0 NET83 NET128 GND GND N18 W=0.92U L=0.18U
MN3 NET68 SN GND GND N18 W=1.86U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.86U L=0.18U
MP1 VDD NET128 NET89 VDD P18 W=3.21U L=0.18U
MP7 VDD NET128 NET77 VDD P18 W=1.68U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET32 NET95 VDD P18 W=0.45U L=0.18U
MP3 VDD SN NET95 VDD P18 W=1.1U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=3.21U L=0.18U
XI9 NET65 NET95 NET32 NET24 TG1G NL=0.19U NW=1.35U PL=0.19U PW=1.35U
.ENDS FFDNSRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSRHD2X                                                           *
* LAST TIME SAVED: DEC  1 15:06:46 2003                                       *
*******************************************************************************
.SUBCKT FFDNSRHD2X Q QN CKN D RN SN
XI32 NET33 NET65 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=1.05U
XI13 NET24 NET32 IVG PW=0.3U NW=0.45U
XI12 QN NET95 IVG PW=2.4U NW=1.6U
XI34 NET128 RN IVG PW=0.81U NW=0.54U
XI10 NET60 NET95 IVG PW=0.84U NW=0.56U
XI5 Q NET60 IVG PW=2.4U NW=1.6U
XI4 NET32 CKN IVG PW=1.2U NW=0.3U
MN1 NET95 NET24 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 SN NET83 GND N18 W=0.58U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN0 NET83 NET128 GND GND N18 W=0.58U L=0.18U
MN3 NET68 SN GND GND N18 W=1.57U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.57U L=0.18U
MP1 VDD NET128 NET89 VDD P18 W=2.2U L=0.18U
MP7 VDD NET128 NET77 VDD P18 W=0.86U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET32 NET95 VDD P18 W=0.45U L=0.18U
MP3 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=2.2U L=0.18U
XI9 NET65 NET95 NET32 NET24 TG1G NW=1.1U PW=1.1U
.ENDS FFDNSRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSRHD1X                                                           *
* LAST TIME SAVED: DEC  1 15:06:23 2003                                       *
*******************************************************************************
.SUBCKT FFDNSRHD1X Q QN CKN D RN SN
XI32 NET33 NET65 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI33 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NET95 IVG PW=1.2U NW=0.8U
XI34 NET128 RN IVG PW=0.64U NW=0.42U
XI10 NET60 NET95 IVG PW=0.64U NW=0.42U
XI5 Q NET60 IVG PW=1.2U NW=0.8U
XI4 NET32 CKN IVG PW=0.78U NW=0.3U
MN1 NET95 NET24 NET62 GND N18 W=0.3U L=0.18U
MN4 NET62 NET60 NET59 GND N18 W=0.3U L=0.18U
MN6 NET95 SN NET83 GND N18 W=0.58U L=0.18U
MN5 NET59 SN GND GND N18 W=0.6U L=0.18U
MN0 NET83 NET128 GND GND N18 W=0.58U L=0.18U
MN3 NET68 SN GND GND N18 W=1.13U L=0.18U
MN2 NET65 NET33 NET68 GND N18 W=1.13U L=0.18U
MP1 VDD NET128 NET89 VDD P18 W=1.6U L=0.18U
MP7 VDD NET128 NET77 VDD P18 W=1U L=0.18U
MP5 NET77 NET60 NET80 VDD P18 W=0.45U L=0.18U
MP4 NET80 NET32 NET95 VDD P18 W=0.45U L=0.18U
MP3 VDD SN NET95 VDD P18 W=0.64U L=0.18U
MP6 NET89 NET33 NET65 VDD P18 W=1.6U L=0.18U
XI9 NET65 NET95 NET32 NET24 TG1G NW=0.7U PW=0.7U
.ENDS FFDNSRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSHDLX                                                            *
* LAST TIME SAVED: DEC  1 15:08:42 2003                                       *
*******************************************************************************
.SUBCKT FFDNSHDLX Q QN CKN D SN
MN1 NET70 NET24 NET38 GND N18 W=0.3U L=0.18U
MN2 NET111 SN GND GND N18 W=0.64U L=0.18U
MN5 NET38 NET36 NET117 GND N18 W=0.3U L=0.18U
MN0 NET117 SN GND GND N18 W=0.6U L=0.18U
MN3 NET62 NET33 NET111 GND N18 W=0.64U L=0.18U
MP7 VDD NET36 NET59 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET70 VDD P18 W=0.64U L=0.18U
MP6 VDD NET33 NET62 VDD P18 W=0.84U L=0.18U
MP4 NET59 NET32 NET70 VDD P18 W=0.45U L=0.18U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI29 NET33 NET62 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET62 NET70 NET32 NET24 TG1G NW=0.5U PW=0.5U
XI12 QN NET70 IVG PW=0.64U NW=0.42U
XI10 NET36 NET70 IVG PW=0.42U NW=0.3U
XI5 Q NET36 IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI4 NET32 CKN IVG PW=0.9U NW=0.3U
.ENDS FFDNSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSHD4X                                                            *
* LAST TIME SAVED: DEC 27 23:13:25 2003                                       *
*******************************************************************************
.SUBCKT FFDNSHD4X Q QN CKN D SN
MN1 NET70 NET24 NET38 GND N18 W=0.3U L=0.18U
MN2 NET111 SN GND GND N18 W=1.86U L=0.18U
MN5 NET38 NET36 NET117 GND N18 W=0.3U L=0.18U
MN0 NET117 SN GND GND N18 W=0.8U L=0.18U
MN3 NET62 NET33 NET111 GND N18 W=1.86U L=0.18U
MP7 VDD NET36 NET59 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET70 VDD P18 W=1.1U L=0.18U
MP6 VDD NET33 NET62 VDD P18 W=2.42U L=0.18U
MP4 NET59 NET32 NET70 VDD P18 W=0.45U L=0.18U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.45U PW=1.62U
XI29 NET33 NET62 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET62 NET70 NET32 NET24 TG1G NL=0.19U NW=1.35U PL=0.19U PW=1.35U
XI12 QN NET70 IVG PW=4.8U NW=3.2U
XI10 NET36 NET70 IVG PW=1.77U NW=1.18U
XI5 Q NET36 IVG PW=4.8U NW=3.2U
XI13 NET24 NET32 IVG PW=0.3U NW=0.48U
XI4 NET32 CKN IVG PW=1.44U NW=0.3U
.ENDS FFDNSHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSHD2X                                                            *
* LAST TIME SAVED: DEC  1 15:08:12 2003                                       *
*******************************************************************************
.SUBCKT FFDNSHD2X Q QN CKN D SN
MN1 NET70 NET24 NET38 GND N18 W=0.3U L=0.18U
MN2 NET111 SN GND GND N18 W=1.57U L=0.18U
MN5 NET38 NET36 NET117 GND N18 W=0.3U L=0.18U
MN0 NET117 SN GND GND N18 W=0.6U L=0.18U
MN3 NET62 NET33 NET111 GND N18 W=1.57U L=0.18U
MP7 VDD NET36 NET59 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET70 VDD P18 W=0.64U L=0.18U
MP6 VDD NET33 NET62 VDD P18 W=1.68U L=0.18U
MP4 NET59 NET32 NET70 VDD P18 W=0.45U L=0.18U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=1.05U
XI29 NET33 NET62 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET62 NET70 NET32 NET24 TG1G NW=1.1U PW=1.1U
XI12 QN NET70 IVG PW=2.4U NW=1.6U
XI10 NET36 NET70 IVG PW=0.84U NW=0.56U
XI5 Q NET36 IVG PW=2.4U NW=1.6U
XI13 NET24 NET32 IVG PW=0.3U NW=0.45U
XI4 NET32 CKN IVG PW=1.2U NW=0.3U
.ENDS FFDNSHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNSHD1X                                                            *
* LAST TIME SAVED: DEC  1 15:07:56 2003                                       *
*******************************************************************************
.SUBCKT FFDNSHD1X Q QN CKN D SN
MN1 NET70 NET24 NET38 GND N18 W=0.3U L=0.18U
MN2 NET111 SN GND GND N18 W=1.13U L=0.18U
MN5 NET38 NET36 NET117 GND N18 W=0.3U L=0.18U
MN0 NET117 SN GND GND N18 W=0.6U L=0.18U
MN3 NET62 NET33 NET111 GND N18 W=1.13U L=0.18U
MP7 VDD NET36 NET59 VDD P18 W=0.45U L=0.18U
MP0 VDD SN NET70 VDD P18 W=0.64U L=0.18U
MP6 VDD NET33 NET62 VDD P18 W=1.22U L=0.18U
MP4 NET59 NET32 NET70 VDD P18 W=0.45U L=0.18U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI29 NET33 NET62 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET62 NET70 NET32 NET24 TG1G NW=0.7U PW=0.7U
XI12 QN NET70 IVG PW=1.2U NW=0.8U
XI10 NET36 NET70 IVG PW=0.64U NW=0.42U
XI5 Q NET36 IVG PW=1.2U NW=0.8U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI4 NET32 CKN IVG PW=0.78U NW=0.3U
.ENDS FFDNSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNRHDLX                                                            *
* LAST TIME SAVED: DEC  1 15:09:40 2003                                       *
*******************************************************************************
.SUBCKT FFDNRHDLX Q QN CKN D RN
MN5 NET36 NET34 GND GND N18 W=0.3U L=0.18U
MN1 NET67 NET24 NET36 GND N18 W=0.3U L=0.18U
MN6 NET67 NET76 GND GND N18 W=0.42U L=0.18U
MN3 NET46 NET33 GND GND N18 W=0.5U L=0.18U
MP1 VDD NET76 NET57 VDD P18 W=1.1U L=0.18U
MP4 NET51 NET32 NET67 VDD P18 W=0.45U L=0.18U
MP7 NET54 NET34 NET51 VDD P18 W=0.45U L=0.18U
MP6 NET57 NET33 NET46 VDD P18 W=1.1U L=0.18U
MP5 VDD NET76 NET54 VDD P18 W=1U L=0.18U
XI29 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI9 NET46 NET67 NET32 NET24 TG1G NW=0.5U PW=0.5U
XI12 QN NET67 IVG PW=0.64U NW=0.42U
XI21 NET76 RN IVG PW=0.64U NW=0.42U
XI5 Q NET34 IVG PW=0.64U NW=0.42U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI10 NET34 NET67 IVG PW=0.42U NW=0.3U
XI4 NET32 CKN IVG PW=0.9U NW=0.3U
.ENDS FFDNRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNRHD4X                                                            *
* LAST TIME SAVED: DEC 27 23:12:08 2003                                       *
*******************************************************************************
.SUBCKT FFDNRHD4X Q QN CKN D RN
MN5 NET36 NET34 GND GND N18 W=0.3U L=0.18U
MN1 NET67 NET24 NET36 GND N18 W=0.3U L=0.18U
MN6 NET67 NET76 GND GND N18 W=0.72U L=0.18U
MN3 NET46 NET33 GND GND N18 W=1.45U L=0.18U
MP1 VDD NET76 NET57 VDD P18 W=3.21U L=0.18U
MP4 NET51 NET32 NET67 VDD P18 W=0.45U L=0.18U
MP7 NET54 NET34 NET51 VDD P18 W=0.45U L=0.18U
MP6 NET57 NET33 NET46 VDD P18 W=3.21U L=0.18U
MP5 VDD NET76 NET54 VDD P18 W=1.68U L=0.18U
XI29 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.45U PW=1.62U
XI9 NET46 NET67 NET32 NET24 TG1G NL=0.19U NW=1.35U PL=0.19U PW=1.35U
XI12 QN NET67 IVG PW=4.8U NW=3.2U
XI21 NET76 RN IVG PW=1.5U NW=1U
XI5 Q NET34 IVG PW=4.8U NW=3.2U
XI13 NET24 NET32 IVG PW=0.3U NW=0.48U
XI10 NET34 NET67 IVG PW=1.77U NW=1.18U
XI4 NET32 CKN IVG PW=1.44U NW=0.3U
.ENDS FFDNRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNRHD2X                                                            *
* LAST TIME SAVED: DEC  1 15:09:12 2003                                       *
*******************************************************************************
.SUBCKT FFDNRHD2X Q QN CKN D RN
MN5 NET36 NET34 GND GND N18 W=0.3U L=0.18U
MN1 NET67 NET24 NET36 GND N18 W=0.3U L=0.18U
MN6 NET67 NET76 GND GND N18 W=0.42U L=0.18U
MN3 NET46 NET33 GND GND N18 W=1.22U L=0.18U
MP1 VDD NET76 NET57 VDD P18 W=2.2U L=0.18U
MP4 NET51 NET32 NET67 VDD P18 W=0.45U L=0.18U
MP7 NET54 NET34 NET51 VDD P18 W=0.45U L=0.18U
MP6 NET57 NET33 NET46 VDD P18 W=2.2U L=0.18U
MP5 VDD NET76 NET54 VDD P18 W=0.86U L=0.18U
XI29 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=1.05U
XI9 NET46 NET67 NET32 NET24 TG1G NW=1.1U PW=1.1U
XI12 QN NET67 IVG PW=2.4U NW=1.6U
XI21 NET76 RN IVG PW=0.81U NW=0.54U
XI5 Q NET34 IVG PW=2.4U NW=1.6U
XI13 NET24 NET32 IVG PW=0.3U NW=0.45U
XI10 NET34 NET67 IVG PW=0.84U NW=0.56U
XI4 NET32 CKN IVG PW=1.2U NW=0.3U
.ENDS FFDNRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNRHD1X                                                            *
* LAST TIME SAVED: DEC  1 15:08:58 2003                                       *
*******************************************************************************
.SUBCKT FFDNRHD1X Q QN CKN D RN
MN5 NET36 NET34 GND GND N18 W=0.3U L=0.18U
MN1 NET67 NET24 NET36 GND N18 W=0.3U L=0.18U
MN6 NET67 NET76 GND GND N18 W=0.42U L=0.18U
MN3 NET46 NET33 GND GND N18 W=0.88U L=0.18U
MP1 VDD NET76 NET57 VDD P18 W=1.6U L=0.18U
MP4 NET51 NET32 NET67 VDD P18 W=0.45U L=0.18U
MP7 NET54 NET34 NET51 VDD P18 W=0.45U L=0.18U
MP6 NET57 NET33 NET46 VDD P18 W=1.6U L=0.18U
MP5 VDD NET76 NET54 VDD P18 W=1U L=0.18U
XI29 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI30 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI9 NET46 NET67 NET32 NET24 TG1G NW=0.7U PW=0.7U
XI12 QN NET67 IVG PW=1.2U NW=0.8U
XI21 NET76 RN IVG PW=0.64U NW=0.42U
XI5 Q NET34 IVG PW=1.2U NW=0.8U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI10 NET34 NET67 IVG PW=0.64U NW=0.42U
XI4 NET32 CKN IVG PW=0.78U NW=0.3U
.ENDS FFDNRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNHDLX                                                             *
* LAST TIME SAVED: DEC  1 15:10:40 2003                                       *
*******************************************************************************
.SUBCKT FFDNHDLX Q QN CKN D
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=0.5U PW=0.5U
XI7 NET46 NET33 IVG PW=0.84U NW=0.5U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NETQ IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.42U NW=0.3U
XI5 Q NETQN IVG PW=0.64U NW=0.42U
XI4 NET32 CKN IVG PW=0.9U NW=0.3U
.ENDS FFDNHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNHD4X                                                             *
* LAST TIME SAVED: DEC  1 15:10:25 2003                                       *
*******************************************************************************
.SUBCKT FFDNHD4X Q QN CKN D
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET24 NET32 TRIIVG NW=0.45U PW=1.62U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=1.35U PW=1.35U
XI7 NET46 NET33 IVG PW=2.42U NW=1.45U
XI13 NET24 NET32 IVG PW=0.3U NW=0.48U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CKN IVG PW=1.44U NW=0.3U
.ENDS FFDNHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNHD2X                                                             *
* LAST TIME SAVED: DEC  1 15:10:10 2003                                       *
*******************************************************************************
.SUBCKT FFDNHD2X Q QN CKN D
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=1.05U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=1.1U PW=1.1U
XI7 NET46 NET33 IVG PW=1.68U NW=1.22U
XI13 NET24 NET32 IVG PW=0.3U NW=0.45U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CKN IVG PW=1.2U NW=0.3U
.ENDS FFDNHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDNHD1X                                                             *
* LAST TIME SAVED: DEC  1 15:09:56 2003                                       *
*******************************************************************************
.SUBCKT FFDNHD1X Q QN CKN D
XI17 NET33 NET46 NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET24 NET32 TRIIVG NW=0.3U PW=0.9U
XI11 NETQ NETQN NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET32 NET24 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=1.22U NW=0.88U
XI13 NET24 NET32 IVG PW=0.3U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CKN IVG PW=0.78U NW=0.3U
.ENDS FFDNHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDHDLX                                                              *
* LAST TIME SAVED: NOV 17 19:14:36 2003                                       *
*******************************************************************************
.SUBCKT FFDHDLX Q QN CK D
XI18 NET33 D NET32 NET24 TRIIVG NW=0.38U PW=0.64U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.5U PW=0.5U
XI7 NET46 NET33 IVG PW=0.84U NW=0.56U
XI13 NET24 NET32 IVG PW=0.42U NW=0.3U
XI20 Q NETQN IVG PW=0.64U NW=0.42U
XI10 NETQN NETQ IVG PW=0.54U NW=0.36U
XI19 QN NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDHD4X                                                              *
* LAST TIME SAVED: DEC  1 15:11:15 2003                                       *
*******************************************************************************
.SUBCKT FFDHD4X Q QN CK D
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI18 NET33 D NET32 NET24 TRIIVG NW=0.78U PW=1.32U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.35U PW=1.35U PL=0.18U NL=0.19U
XI7 NET46 NET33 IVG PW=2.52U NW=1.68U
XI13 NET24 NET32 IVG PW=0.93U NW=0.3U
XI12 QN NETQ IVG PW=4.8U NW=3.2U
XI10 NETQN NETQ IVG PW=1.77U NW=1.18U
XI5 Q NETQN IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=0.3U NW=0.8U
.ENDS FFDHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDHD2XSPG                                                           *
* LAST TIME SAVED: NOV 17 15:15:23 2003                                       *
*******************************************************************************
.SUBCKT FFDHD2XSPG Q QN CK D
XI18 NET33 D NET32 NET24 TRIIVG NW=0.54U PW=0.96U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFDHD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDHD2X                                                              *
* LAST TIME SAVED: NOV 17 15:14:00 2003                                       *
*******************************************************************************
.SUBCKT FFDHD2X Q QN CK D
XI18 NET33 D NET32 NET24 TRIIVG NW=0.54U PW=0.96U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=1.1U PW=1.1U
XI7 NET46 NET33 IVG PW=1.72U NW=1.22U
XI13 NET24 NET32 IVG PW=0.69U NW=0.3U
XI12 QN NETQ IVG PW=2.4U NW=1.6U
XI10 NETQN NETQ IVG PW=0.84U NW=0.56U
XI5 Q NETQN IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=0.3U NW=0.45U
.ENDS FFDHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDHD1X                                                              *
* LAST TIME SAVED: NOV 17 14:53:51 2003                                       *
*******************************************************************************
.SUBCKT FFDHD1X Q QN CK D
XI18 NET33 D NET32 NET24 TRIIVG NW=0.42U PW=0.84U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQ NETQN NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI9 NET46 NETQ NET24 NET32 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQ IVG PW=1.2U NW=0.8U
XI10 NETQN NETQ IVG PW=0.64U NW=0.42U
XI5 Q NETQN IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.3U NW=0.3U
.ENDS FFDHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDCRHDLX                                                            *
* LAST TIME SAVED: MAR  4 14:28:38 2003                                       *
*******************************************************************************
.SUBCKT FFDCRHDLX Q QN CK D RN
XI18 NET63 RN D ND2G PW=0.6U NW=0.5U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=0.93U NW=0.62U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=0.64U NW=0.42U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=0.64U NW=0.42U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFDCRHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDCRHD4X                                                            *
* LAST TIME SAVED: MAR  4 14:28:06 2003                                       *
*******************************************************************************
.SUBCKT FFDCRHD4X Q QN CK D RN
XI18 NET63 RN D ND2G PW=1.47U NW=1.18U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.6U PW=0.6U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.18U PW=1.18U
XI7 NET46 NET33 IVG PW=3.44U NW=2.3U
XI13 NET24 NET32 IVG PW=0.96U NW=0.48U
XI12 QN NETQN IVG PW=4.8U NW=3.2U
XI10 NETQ NETQN IVG PW=1.68U NW=1.14U
XI5 Q NETQ IVG PW=4.8U NW=3.2U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFDCRHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDCRHD2X                                                            *
* LAST TIME SAVED: MAR  4 14:27:38 2003                                       *
*******************************************************************************
.SUBCKT FFDCRHD2X Q QN CK D RN
XI18 NET63 RN D ND2G PW=0.96U NW=0.8U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI6 NET63 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=1.1U PW=1.1U
XI7 NET46 NET33 IVG PW=1.72U NW=1.18U
XI13 NET24 NET32 IVG PW=0.84U NW=0.42U
XI12 QN NETQN IVG PW=2.4U NW=1.6U
XI10 NETQ NETQN IVG PW=0.84U NW=0.56U
XI5 Q NETQ IVG PW=2.4U NW=1.6U
XI4 NET32 CK IVG PW=1.2U NW=0.6U
.ENDS FFDCRHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FFDCRHD1X                                                            *
* LAST TIME SAVED: MAR  4 14:27:07 2003                                       *
*******************************************************************************
.SUBCKT FFDCRHD1X Q QN CK D RN
XI18 NET34 RN D ND2G PW=0.66U NW=0.55U
XI17 NET33 NET46 NET24 NET32 TRIIVG NW=0.3U PW=0.42U
XI11 NETQN NETQ NET32 NET24 TRIIVG NW=0.3U PW=0.42U
XI6 NET34 NET33 NET32 NET24 TG1G NW=0.42U PW=0.42U
XI9 NET46 NETQN NET24 NET32 TG1G NW=0.7U PW=0.7U
XI7 NET46 NET33 IVG PW=1.28U NW=0.86U
XI13 NET24 NET32 IVG PW=0.6U NW=0.3U
XI12 QN NETQN IVG PW=1.2U NW=0.8U
XI10 NETQ NETQN IVG PW=0.64U NW=0.42U
XI5 Q NETQ IVG PW=1.2U NW=0.8U
XI4 NET32 CK IVG PW=0.84U NW=0.42U
.ENDS FFDCRHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHHDLX                                                              *
* LAST TIME SAVED: AUG 30 10:29:35 2002                                       *
*******************************************************************************
.SUBCKT FAHHDLX CO S A B CI
XI21 NET132 NET105 NET117 NET123 TG1G NW=0.6U PW=0.6U
XI20 NET138 NET123 B NET132 TG1G NW=0.8U PW=0.8U
XI18 NET138 NET117 NET132 B TG1G NW=0.8U PW=0.8U
XI17 NET124 NET111 NET123 NET117 TG1G NW=0.6U PW=0.6U
XI14 NET130 NET111 NET117 NET123 TG1G NW=0.6U PW=0.6U
XI12 NET130 NET105 NET123 NET117 TG1G NW=0.6U PW=0.6U
XI6 NET_92 NET123 NET132 B TG1G NW=0.8U PW=0.8U
XI4 NET_92 NET117 B NET132 TG1G NW=0.8U PW=0.8U
XI15 S NET111 IVG PW=0.64U NW=0.42U
XI13 CO NET105 IVG PW=0.64U NW=0.42U
XI26 NET124 NET130 IVG PW=0.45U NW=0.3U
XI22 NET138 A IVG PW=0.9U NW=0.6U
XI25 NET130 CI IVG PW=0.45U NW=0.3U
XI24 NET132 B IVG PW=0.45U NW=0.3U
XI23 NET_92 NET138 IVG PW=0.45U NW=0.3U
.ENDS FAHHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHHD4X                                                              *
* LAST TIME SAVED: AUG 30 10:29:33 2002                                       *
*******************************************************************************
.SUBCKT FAHHD4X CO S A B CI
XI11 NET_121 NET130 IVG PW=1.8U NW=1.2U
XI10 NET132 B IVG PW=3U NW=2U
XI7 NET130 CI IVG PW=2.4U NW=1.6U
XI3 NET_113 NET138 IVG PW=3.0U NW=2.0U
XI2 NET138 A IVG PW=3.44U NW=2.44U
XI15 S NET111 IVG PW=4.8U NW=3.2U
XI13 CO NET105 IVG PW=4.8U NW=3.2U
XI18 NET138 NET_135 NET132 B TG1G NW=2.0U PW=2.0U
XI20 NET138 NET_134 B NET132 TG1G NW=2.0U PW=2.0U
XI1 NET130 NET105 NET_134 NET_135 TG1G NW=1.18U PW=1.2U
XI0 NET130 NET111 NET_135 NET_134 TG1G NW=1.18U PW=1.2U
XI6 NET_113 NET_134 NET132 B TG1G NW=2.0U PW=2.0U
XI4 NET_113 NET_135 B NET132 TG1G NW=2.0U PW=2.0U
XI17 NET_121 NET111 NET_134 NET_135 TG1G NW=1.18U PW=1.2U
XI5 NET132 NET105 NET_135 NET_134 TG1G NW=1.18U PW=1.2U
.ENDS FAHHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHHD2X                                                              *
* LAST TIME SAVED: AUG 30 10:29:30 2002                                       *
*******************************************************************************
.SUBCKT FAHHD2X CO S A B CI
XI2 NET138 A IVG PW=3.44U NW=2.44U
XI3 NET_9 NET138 IVG PW=3.0U NW=2.0U
XI7 NET130 CI IVG PW=2.4U NW=1.6U
XI10 NET132 B IVG PW=3U NW=2U
XI11 NET_17 NET130 IVG PW=1.8U NW=1.2U
XI13 CO NET105 IVG PW=2.4U NW=1.6U
XI15 S NET111 IVG PW=2.4U NW=1.6U
XI4 NET_9 NET_51 B NET132 TG1G NW=2.0U PW=2.0U
XI6 NET_9 NET_50 NET132 B TG1G NW=2.0U PW=2.0U
XI12 NET130 NET105 NET_50 NET_51 TG1G NW=1.18U PW=1.2U
XI8 NET130 NET111 NET_51 NET_50 TG1G NW=1.18U PW=1.2U
XI17 NET_17 NET111 NET_50 NET_51 TG1G NW=1.18U PW=1.2U
XI18 NET138 NET_51 NET132 B TG1G NW=2.0U PW=2.0U
XI20 NET138 NET_50 B NET132 TG1G NW=2.0U PW=2.0U
XI14 NET132 NET105 NET_51 NET_50 TG1G NW=1.18U PW=1.2U
.ENDS FAHHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHHD1X                                                              *
* LAST TIME SAVED: AUG 30 10:29:25 2002                                       *
*******************************************************************************
.SUBCKT FAHHD1X CO S A B CI
XI22 NET130 NET111 NET117 NET123 TG1G NW=0.8U PW=0.8U
XI31 NET_92 NET117 B NET132 TG1G NW=0.9U PW=1.3U
XI18 NET138 NET117 NET132 B TG1G NW=0.9U PW=1.3U
XI17 NET_68 NET111 NET123 NET117 TG1G NW=0.8U PW=0.8U
XI24 NET132 NET105 NET117 NET123 TG1G NW=0.8U PW=0.8U
XI23 NET130 NET105 NET123 NET117 TG1G NW=0.8U PW=0.8U
XI32 NET_92 NET123 NET132 B TG1G NW=0.9U PW=1.3U
XI33 NET138 NET123 B NET132 TG1G NW=0.9U PW=1.3U
XI15 S NET111 IVG PW=1.2U NW=0.8U
XI13 CO NET105 IVG PW=1.2U NW=0.8U
XI11 NET_68 NET130 IVG PW=0.9U NW=0.6U
XI10 NET132 B IVG PW=1.4U NW=1.0U
XI7 NET130 CI IVG PW=1.2U NW=0.8U
XI3 NET_92 NET138 IVG PW=1.65U NW=1.12U
XI2 NET138 A IVG PW=1.72U NW=1.22U
.ENDS FAHHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHDLX                                                               *
* LAST TIME SAVED: AUG 30 10:29:42 2002                                       *
*******************************************************************************
.SUBCKT FAHDLX CO S A B CI
XI5 CO NET28 IVG PW=0.64U NW=0.42U
XI9 NET9 NET15 IVG PW=0.9U NW=0.6U
XI2 NET11 CI IVG PW=0.64U NW=0.42U
XI10 NET13 A IVG PW=0.9U NW=0.6U
XI1 NET15 B IVG PW=0.9U NW=0.6U
XI8 S NET32 IVG PW=0.64U NW=0.42U
XI4 NET13 NET52 NET9 NET15 TG1G NW=0.6U PW=0.6U
XI0 NET13 NET44 NET15 NET9 TG1G NW=0.6U PW=0.6U
XI3 NET11 NET28 NET52 NET44 TG1G NW=0.6U PW=0.6U
XI7 NET52 NET32 CI NET11 TG1G NW=0.6U PW=0.6U
XI12 NET15 NET28 NET44 NET52 TG1G NW=0.6U PW=0.6U
XI6 NET44 NET32 NET11 CI TG1G NW=0.6U PW=0.6U
MP1 NET44 NET13 NET15 GND N18 W=0.64U L=0.18U
MN1 NET52 NET13 NET9 GND N18 W=0.64U L=0.18U
MP0 NET9 NET13 NET44 VDD P18 W=0.96U L=0.18U
MP2 NET15 NET13 NET52 VDD P18 W=0.96U L=0.18U
.ENDS FAHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHD4X                                                               *
* LAST TIME SAVED: DEC 27 23:29:18 2003                                       *
*******************************************************************************
.SUBCKT FAHD4X CO S A B CI
MP2 NET45 NET47 NET7 VDD P18 W=1.5U L=0.18U
MP0 NET51 NET47 NET17 VDD P18 W=1.2U L=0.18U
MN1 NET7 NET47 NET51 GND N18 W=1.0U L=0.18U
MP1 NET17 NET47 NET45 GND N18 W=1.0U L=0.18U
XI6 NET17 NET28 NET49 CI TG1G NW=1.2U PW=1.2U
XI12 NET45 NET32 NET17 NET7 TG1G NW=1.0U PW=1.0U
XI7 NET7 NET28 CI NET49 TG1G NL=0.19U NW=1.2U PL=0.19U PW=1.2U
XI3 NET49 NET32 NET7 NET17 TG1G NW=1.0U PW=1.0U
XI0 NET47 NET17 NET45 NET51 TG1G NL=0.19U NW=1.2U PL=0.19U PW=1.2U
XI4 NET47 NET7 NET51 NET45 TG1G NL=0.19U NW=1.2U PL=0.19U PW=1.2U
XI10 NET47 A IVG PW=1.72U NW=1.2U
XI8 S NET28 IVG PW=4.8U NW=3.2U
XI1 NET45 B IVG PW=1.72U NW=1.2U
XI2 NET49 CI IVG PL=0.19U PW=1.4U NW=1.0U
XI9 NET51 NET45 IVG PW=1.72U NW=1.2U
XI5 CO NET32 IVG PW=4.8U NW=3.2U
.ENDS FAHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHD2X                                                               *
* LAST TIME SAVED: DEC 27 23:30:33 2003                                       *
*******************************************************************************
.SUBCKT FAHD2X CO S A B CI
XI10 NET13 A IVG PW=1.72U NW=1.2U
XI5 CO NET28 IVG PW=2.4U NW=1.6U
XI8 S NET32 IVG PW=2.4U NW=1.6U
XI16 NET9 NET15 IVG PW=1.72U NW=1.2U
XI15 NET15 B IVG PW=1.72U NW=1.2U
XI2 NET11 CI IVG PW=1.2U NW=0.8U PL=0.19U NL=0.18U
XI11 NET13 NET52 NET9 NET15 TG1G NW=1.0U PW=1.0U
XI14 NET52 NET32 CI NET11 TG1G NW=1.0U PW=1.0U
XI12 NET15 NET28 NET44 NET52 TG1G NW=0.8U PW=0.8U
XI3 NET11 NET28 NET52 NET44 TG1G NW=0.8U PW=0.8U
XI0 NET13 NET44 NET15 NET9 TG1G NW=1.0U PW=1.0U
XI13 NET44 NET32 NET11 CI TG1G NW=1.0U PW=1.0U
MN1 NET52 NET13 NET9 GND N18 W=1.0U L=0.18U
MN0 NET44 NET13 NET15 GND N18 W=1.0U L=0.18U
MP1 NET15 NET13 NET52 VDD P18 W=1.5U L=0.18U
MP0 NET9 NET13 NET44 VDD P18 W=1.5U L=0.19U
.ENDS FAHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FAHD1X                                                               *
* LAST TIME SAVED: AUG 30 10:29:37 2002                                       *
*******************************************************************************
.SUBCKT FAHD1X CO S A B CI
MP2 NET117 NET119 NET_103 VDD P18 W=1.2U L=0.18U
MP0 NET109 NET119 NET_102 VDD P18 W=1.2U L=0.18U
MP1 NET_102 NET119 NET117 GND N18 W=0.8U L=0.18U
MN1 NET_103 NET119 NET109 GND N18 W=0.8U L=0.18U
XI12 NET117 NET_6 NET_102 NET_103 TG1G NW=0.6U PW=0.6U
XI13 NET119 NET_103 NET109 NET117 TG1G NW=0.8U PW=0.8U
XI18 NET115 NET_6 NET_103 NET_102 TG1G NW=0.6U PW=0.6U
XI14 NET_102 NET108 NET115 CI TG1G NW=0.8U PW=0.8U
XI0 NET119 NET_102 NET117 NET109 TG1G NW=0.8U PW=0.8U
XI15 NET_103 NET108 CI NET115 TG1G NW=0.8U PW=0.8U
XI16 NET109 NET117 IVG PW=1.72U NW=1.2U
XI8 S NET108 IVG PW=1.2U NW=0.8U
XI5 CO NET_6 IVG PW=1.2U NW=0.8U
XI2 NET115 CI IVG PW=0.9U NW=0.6U
XI1 NET117 B IVG PW=1.72U NW=1.2U
XI17 NET119 A IVG PW=1.72U NW=1.2U
.ENDS FAHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IVGII                                                                *
* LAST TIME SAVED: SEP 10 14:37:23 2001                                       *
*******************************************************************************
.SUBCKT IVGII Z A PL=0.18U PW=0.24U NL=0.18U NW=0.24U
MN0 Z A GND GND N18 W=NW L=NL
MP0 VDD A Z VDD P18 W=PW L=PL
.ENDS IVGII


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL4HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:32:51 2002                                       *
*******************************************************************************
.SUBCKT DEL4HD2X Z A
XI4 Z NET23 IVGII PL=0.18U PW=2.4U NL=0.18U NW=1.6U
XI5 NET23 NET21 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI6 NET21 NET19 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI7 NET19 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL4HD1XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:32:51 2002                                       *
*******************************************************************************
.SUBCKT DEL4HD1XSPG Z A
XI0 Z NET6 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI1 NET6 NET8 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL4HD1XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL4HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:32:49 2002                                       *
*******************************************************************************
.SUBCKT DEL4HD1X Z A
XI0 Z NET6 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI1 NET6 NET8 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.72U PW=0.45U NL=0.72U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL3HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:32:47 2002                                       *
*******************************************************************************
.SUBCKT DEL3HD2X Z A
XI0 Z NET6 IVGII PL=0.18U PW=2.4U NL=0.18U NW=1.6U
XI1 NET6 NET8 IVGII PL=0.54U PW=0.45U NL=0.54U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.54U PW=0.45U NL=0.54U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL3HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:32:46 2002                                       *
*******************************************************************************
.SUBCKT DEL3HD1X Z A
XI0 Z NET6 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI1 NET6 NET8 IVGII PL=0.54U PW=0.45U NL=0.54U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.54U PW=0.45U NL=0.54U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL3HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL2HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:32:44 2002                                       *
*******************************************************************************
.SUBCKT DEL2HD2X Z A
XI7 NET19 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI4 Z NET23 IVGII PL=0.18U PW=2.4U NL=0.18U NW=1.6U
XI5 NET23 NET21 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
XI6 NET21 NET19 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
.ENDS DEL2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL2HD1XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:32:42 2002                                       *
*******************************************************************************
.SUBCKT DEL2HD1XSPG Z A
XI4 Z NET13 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI5 NET13 NET11 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
XI6 NET11 NET9 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
XI7 NET9 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL2HD1XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL2HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:32:41 2002                                       *
*******************************************************************************
.SUBCKT DEL2HD1X Z A
XI0 Z NET6 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI1 NET6 NET8 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.36U PW=0.45U NL=0.36U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL1HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:32:39 2002                                       *
*******************************************************************************
.SUBCKT DEL1HD2X Z A
XI0 Z NET6 IVGII PL=0.18U PW=2.4U NL=0.18U NW=1.6U
XI1 NET6 NET8 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI2 NET8 NET10 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI3 NET10 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL1HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL1HD1XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:32:37 2002                                       *
*******************************************************************************
.SUBCKT DEL1HD1XSPG Z A
XI4 Z NET13 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
XI5 NET13 NET11 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI6 NET11 NET9 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI7 NET9 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
.ENDS DEL1HD1XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DEL1HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:32:35 2002                                       *
*******************************************************************************
.SUBCKT DEL1HD1X Z A
XI3 NET4 A IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI2 NET6 NET4 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI1 NET8 NET6 IVGII PL=0.18U PW=0.45U NL=0.18U NW=0.3U
XI0 Z NET8 IVGII PL=0.18U PW=1.2U NL=0.18U NW=0.8U
.ENDS DEL1HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHDLX                                                            *
* LAST TIME SAVED: AUG 30 10:44:38 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHDLX Z A E
MN2 NET9 NET27 GND GND N18 W=0.42U L=0.18U
MN1 NET9 A GND GND N18 W=0.42U L=0.18U
MN0 Z NET9 GND GND N18 W=0.42U L=0.18U
MP4 VDD NET14 Z VDD P18 W=0.64U L=0.18U
MP1 VDD E NET14 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET14 VDD P18 W=0.64U L=0.18U
XI6 NET9 NET14 E NET27 TG1G NW=0.42U PW=0.42U
XI3 NET27 E IVG PW=0.42U NW=0.30U
.ENDS BUFTSHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD8X                                                            *
* LAST TIME SAVED: AUG 30 10:44:36 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD8X Z A E
XI3 NET5 E IVG PW=0.48U NW=0.32U
XI6 NET24 NET17 E NET5 TG1G NW=1.2U PW=1.72U
MP4 VDD NET17 Z VDD P18 W=9.6U L=0.18U
MP1 VDD E NET17 VDD P18 W=1.2U L=0.18U
MP0 VDD A NET17 VDD P18 W=3.44U L=0.18U
MN2 NET24 NET5 GND GND N18 W=0.8U L=0.18U
MN1 NET24 A GND GND N18 W=2.4U L=0.18U
MN0 Z NET24 GND GND N18 W=6.4U L=0.18U
.ENDS BUFTSHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD3X                                                            *
* LAST TIME SAVED: AUG 30 10:44:24 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD3X Z A E
XI3 NET5 E IVG PW=0.45U NW=0.30U
XI6 NET24 NET17 E NET5 TG1G NW=0.6U PW=0.6U
MP4 VDD NET17 Z VDD P18 W=3.6U L=0.18U
MP1 VDD E NET17 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET17 VDD P18 W=1.44U L=0.18U
MN2 NET24 NET5 GND GND N18 W=0.42U L=0.18U
MN1 NET24 A GND GND N18 W=0.96U L=0.18U
MN0 Z NET24 GND GND N18 W=2.4U L=0.18U
.ENDS BUFTSHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD20X                                                           *
* LAST TIME SAVED: AUG 30 10:44:20 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD20X Z A E
MN0 Z NET9 GND GND N18 W=16U L=0.18U
MN1 NET9 A GND GND N18 W=5.6U L=0.18U
MN2 NET9 NET27 GND GND N18 W=2.0U L=0.18U
MP0 VDD A NET14 VDD P18 W=8.4U L=0.18U
MP1 VDD E NET14 VDD P18 W=2.84U L=0.18U
MP4 VDD NET14 Z VDD P18 W=24U L=0.18U
XI6 NET9 NET14 E NET27 TG1G NW=3.5U PW=3.5U
XI3 NET27 E IVG PW=1.2U NW=0.8U
.ENDS BUFTSHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD1X                                                            *
* LAST TIME SAVED: AUG 30 10:44:08 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD1X Z A E
XI3 NET9 E IVG PW=0.45U NW=0.30U
XI6 NET24 NET17 E NET9 TG1G NW=0.4U PW=0.4U
MP4 VDD NET17 Z VDD P18 W=1.2U L=0.18U
MP1 VDD E NET17 VDD P18 W=0.6U L=0.18U
MP0 VDD A NET17 VDD P18 W=0.64U L=0.18U
MN2 NET24 NET9 GND GND N18 W=0.42U L=0.18U
MN1 NET24 A GND GND N18 W=0.42U L=0.18U
MN0 Z NET24 GND GND N18 W=0.8U L=0.18U
.ENDS BUFTSHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD16X                                                           *
* LAST TIME SAVED: AUG 30 10:44:12 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD16X Z A E
XI3 NET5 E IVG PW=0.96U NW=0.64U
XI6 NET24 NET17 E NET5 TG1G NW=2.36U PW=2.36U
MP4 VDD NET17 Z VDD P18 W=19.2U L=0.18U
MP1 VDD E NET17 VDD P18 W=2.4U L=0.18U
MP0 VDD A NET17 VDD P18 W=6.88U L=0.18U
MN2 NET24 NET5 GND GND N18 W=1.6U L=0.18U
MN1 NET24 A GND GND N18 W=4.8U L=0.18U
MN0 Z NET24 GND GND N18 W=12.8U L=0.18U
.ENDS BUFTSHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFTSHD12X                                                           *
* LAST TIME SAVED: AUG 30 10:44:10 2002                                       *
*******************************************************************************
.SUBCKT BUFTSHD12X Z A E
MN0 Z NET9 GND GND N18 W=9.6U L=0.18U
MN1 NET9 A GND GND N18 W=3.2U L=0.18U
MN2 NET9 NET27 GND GND N18 W=1.2U L=0.18U
MP0 VDD A NET14 VDD P18 W=4.8U L=0.18U
MP1 VDD E NET14 VDD P18 W=1.72U L=0.18U
MP4 VDD NET14 Z VDD P18 W=14.4U L=0.18U
XI6 NET9 NET14 E NET27 TG1G NW=1.8U PW=1.8U
XI3 NET27 E IVG PW=0.72U NW=0.48U
.ENDS BUFTSHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHDLX                                                              *
* LAST TIME SAVED: AUG 30 10:31:47 2002                                       *
*******************************************************************************
.SUBCKT BUFHDLX Z A
XI0 NET4 A IVG PW=0.6U NW=0.42U
XI1 Z NET4 IVG PW=0.6U NW=0.42U
.ENDS BUFHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD8XSPG                                                           *
* LAST TIME SAVED: AUG 30 10:31:45 2002                                       *
*******************************************************************************
.SUBCKT BUFHD8XSPG Z A
XI0 NET4 A IVG PW=3U NW=2U
XI1 Z NET4 IVG PW=9.6U NW=6.4U
.ENDS BUFHD8XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD8X                                                              *
* LAST TIME SAVED: AUG 30 10:31:44 2002                                       *
*******************************************************************************
.SUBCKT BUFHD8X Z A
XI0 NET4 A IVG PW=3U NW=2U
XI1 Z NET4 IVG PW=9.6U NW=6.4U
.ENDS BUFHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD4X                                                              *
* LAST TIME SAVED: AUG 30 10:31:42 2002                                       *
*******************************************************************************
.SUBCKT BUFHD4X Z A
XI1 Z NET6 IVG PW=4.8U NW=3.2U
XI0 NET6 A IVG PW=1.68U NW=1.18U
.ENDS BUFHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD3X                                                              *
* LAST TIME SAVED: AUG 30 10:31:40 2002                                       *
*******************************************************************************
.SUBCKT BUFHD3X Z A
XI0 NET4 A IVG PW=1.2U NW=0.8U
XI1 Z NET4 IVG PW=3.6U NW=2.4U
.ENDS BUFHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD2X                                                              *
* LAST TIME SAVED: AUG 30 10:31:37 2002                                       *
*******************************************************************************
.SUBCKT BUFHD2X Z A
XI1 Z NET6 IVG PW=2.4U NW=1.6U
XI0 NET6 A IVG PW=0.9U NW=0.6U
.ENDS BUFHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD20X                                                             *
* LAST TIME SAVED: AUG 30 10:31:38 2002                                       *
*******************************************************************************
.SUBCKT BUFHD20X Z A
XI1 Z NET6 IVG PW=24U NW=16U
XI0 NET6 A IVG PW=6U NW=4U
.ENDS BUFHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD1X                                                              *
* LAST TIME SAVED: AUG 30 10:31:32 2002                                       *
*******************************************************************************
.SUBCKT BUFHD1X Z A
XI0 NET4 A IVG PW=0.64U NW=0.42U
XI1 Z NET4 IVG PW=1.2U NW=0.8U
.ENDS BUFHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD16X                                                             *
* LAST TIME SAVED: AUG 30 10:31:35 2002                                       *
*******************************************************************************
.SUBCKT BUFHD16X Z A
XI1 Z NET6 IVG PW=19.2U NW=12.8U
XI0 NET6 A IVG PW=4.8U NW=3.2U
.ENDS BUFHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFHD12X                                                             *
* LAST TIME SAVED: AUG 30 10:31:34 2002                                       *
*******************************************************************************
.SUBCKT BUFHD12X Z A
XI1 Z NET6 IVG PW=14.4U NW=9.6U
XI0 NET6 A IVG PW=3.4U NW=2.4U
.ENDS BUFHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHDLX                                                           *
* LAST TIME SAVED: AUG 30 10:32:08 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHDLX Z A
XI0 NET4 A IVG PW=0.45U NW=0.3U
XI1 Z NET4 IVG PW=0.74U NW=0.3U
.ENDS BUFCLKHDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD8X                                                           *
* LAST TIME SAVED: AUG 30 10:32:04 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD8X Z A
XI0 NET4 A IVG PW=2.4U NW=1.2U
XI1 Z NET4 IVG PW=9.6U NW=4.4U
.ENDS BUFCLKHD8X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD80X                                                          *
* LAST TIME SAVED: AUG 30 10:32:05 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD80X Z A
XI1 Z NET6 IVG PW=96U NW=42U
XI0 NET6 A IVG PW=14.4U NW=7.2U
.ENDS BUFCLKHD80X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD4X                                                           *
* LAST TIME SAVED: AUG 30 10:32:00 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD4X Z A
XI1 Z NET6 IVG PW=4.8U NW=2.2U
XI0 NET6 A IVG PW=1.2U NW=0.6U
.ENDS BUFCLKHD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD40X                                                          *
* LAST TIME SAVED: AUG 30 10:32:02 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD40X Z A
XI0 NET4 A IVG PW=8U NW=3.8U
XI1 Z NET4 IVG PW=48U NW=20U
.ENDS BUFCLKHD40X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD3X                                                           *
* LAST TIME SAVED: AUG 30 10:31:56 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD3X Z A
XI0 NET4 A IVG PW=1U NW=0.5U
XI1 Z NET4 IVG PW=3.6U NW=1.6U
.ENDS BUFCLKHD3X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD30X                                                          *
* LAST TIME SAVED: AUG 30 10:31:59 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD30X Z A
XI1 Z NET6 IVG PW=36U NW=16U
XI0 NET6 A IVG PW=5.6U NW=2.8U
.ENDS BUFCLKHD30X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD2X                                                           *
* LAST TIME SAVED: AUG 30 10:31:53 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD2X Z A
XI1 Z NET6 IVG PW=2.4U NW=1.1U
XI0 NET6 A IVG PW=1.2U NW=0.6U
.ENDS BUFCLKHD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD20X                                                          *
* LAST TIME SAVED: AUG 30 10:31:55 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD20X Z A
XI1 Z NET6 IVG PW=24U NW=11U
XI0 NET6 A IVG PW=4.2U NW=2.2U
.ENDS BUFCLKHD20X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD1X                                                           *
* LAST TIME SAVED: AUG 30 10:31:48 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD1X Z A
XI0 NET4 A IVG PW=0.9U NW=0.42U
XI1 Z NET4 IVG PW=1.2U NW=0.5U
.ENDS BUFCLKHD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD16X                                                          *
* LAST TIME SAVED: AUG 30 10:31:51 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD16X Z A
XI1 Z NET6 IVG PW=19.2U NW=8.4U
XI0 NET6 A IVG PW=4U NW=2U
.ENDS BUFCLKHD16X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BUFCLKHD12X                                                          *
* LAST TIME SAVED: AUG 30 10:31:50 2002                                       *
*******************************************************************************
.SUBCKT BUFCLKHD12X Z A
XI1 Z NET6 IVG PW=14.4U NW=6.4U
XI0 NET6 A IVG PW=3.44U NW=1.48U
.ENDS BUFCLKHD12X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI33HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:31:30 2002                                       *
*******************************************************************************
.SUBCKT AOI33HDLX Z A B C D E F
MP5 NET8 E Z VDD P18 W=0.84U L=0.18U
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP4 NET8 D Z VDD P18 W=0.84U L=0.18U
MP2 NET8 F Z VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN7 NET55 D GND GND N18 W=0.58U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN6 NET45 E NET55 GND N18 W=0.58U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 Z C NET12 GND N18 W=0.58U L=0.18U
MN0 Z F NET45 GND N18 W=0.58U L=0.18U
.ENDS AOI33HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI33HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:31:29 2002                                       *
*******************************************************************************
.SUBCKT AOI33HD4X Z A B C D E F
XI4 NET35 NET46 IVG PW=1.6U NW=1.06U
XI5 Z NET35 IVG PW=4.8U NW=3.2U
MP5 NET8 E NET46 VDD P18 W=0.84U L=0.18U
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP4 NET8 D NET46 VDD P18 W=0.84U L=0.18U
MP2 NET8 F NET46 VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN7 NET55 D GND GND N18 W=0.58U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN6 NET45 E NET55 GND N18 W=0.58U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 NET46 C NET12 GND N18 W=0.58U L=0.18U
MN0 NET46 F NET45 GND N18 W=0.58U L=0.18U
.ENDS AOI33HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI33HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:31:27 2002                                       *
*******************************************************************************
.SUBCKT AOI33HD2X Z A B C D E F
MP5 NET8 E Z VDD P18 W=3.2U L=0.18U
MP3 VDD B NET8 VDD P18 W=3.2U L=0.18U
MP4 NET8 D Z VDD P18 W=3.2U L=0.18U
MP2 NET8 F Z VDD P18 W=3.2U L=0.18U
MP1 VDD C NET8 VDD P18 W=3.2U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.2U L=0.18U
MN7 NET55 D GND GND N18 W=2.2U L=0.18U
MN5 NET37 A GND GND N18 W=2.2U L=0.18U
MN6 NET45 E NET55 GND N18 W=2.2U L=0.18U
MN4 NET12 B NET37 GND N18 W=2.2U L=0.18U
MN1 Z C NET12 GND N18 W=2.2U L=0.18U
MN0 Z F NET45 GND N18 W=2.2U L=0.18U
.ENDS AOI33HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI33HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:31:26 2002                                       *
*******************************************************************************
.SUBCKT AOI33HD1X Z A B C D E F
MP5 NET8 E Z VDD P18 W=1.6U L=0.18U
MP3 VDD B NET8 VDD P18 W=1.6U L=0.18U
MP4 NET8 D Z VDD P18 W=1.6U L=0.18U
MP2 NET8 F Z VDD P18 W=1.6U L=0.18U
MP1 VDD C NET8 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.6U L=0.18U
MN7 NET55 D GND GND N18 W=1.1U L=0.18U
MN5 NET37 A GND GND N18 W=1.1U L=0.18U
MN6 NET45 E NET55 GND N18 W=1.1U L=0.18U
MN4 NET12 B NET37 GND N18 W=1.1U L=0.18U
MN1 Z C NET12 GND N18 W=1.1U L=0.18U
MN0 Z F NET45 GND N18 W=1.1U L=0.18U
.ENDS AOI33HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI32HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:31:22 2002                                       *
*******************************************************************************
.SUBCKT AOI32HDLX Z A B C D E
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP4 NET8 D Z VDD P18 W=0.84U L=0.18U
MP2 NET8 E Z VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN6 NET45 D GND GND N18 W=0.52U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 Z C NET12 GND N18 W=0.58U L=0.18U
MN0 Z E NET45 GND N18 W=0.52U L=0.18U
.ENDS AOI32HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI32HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:31:22 2002                                       *
*******************************************************************************
.SUBCKT AOI32HD4X Z A B C D E
XI4 NET69 NET42 IVG PW=1.6U NW=1.06U
XI5 Z NET69 IVG PW=4.8U NW=3.2U
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP4 NET8 D NET42 VDD P18 W=0.84U L=0.18U
MP2 NET8 E NET42 VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN6 NET45 D GND GND N18 W=0.52U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 NET42 C NET12 GND N18 W=0.58U L=0.18U
MN0 NET42 E NET45 GND N18 W=0.52U L=0.18U
.ENDS AOI32HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI32HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:31:19 2002                                       *
*******************************************************************************
.SUBCKT AOI32HD2X Z A B C D E
MP3 VDD B NET8 VDD P18 W=3.2U L=0.18U
MP4 NET8 D Z VDD P18 W=3.2U L=0.18U
MP2 NET8 E Z VDD P18 W=3.2U L=0.18U
MP1 VDD C NET8 VDD P18 W=3.2U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.2U L=0.18U
MN5 NET37 A GND GND N18 W=2.2U L=0.18U
MN6 NET45 D GND GND N18 W=2.0U L=0.18U
MN4 NET12 B NET37 GND N18 W=2.2U L=0.18U
MN1 Z C NET12 GND N18 W=2.2U L=0.18U
MN0 Z E NET45 GND N18 W=2.0U L=0.18U
.ENDS AOI32HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI32HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:31:18 2002                                       *
*******************************************************************************
.SUBCKT AOI32HD1X Z A B C D E
MP3 VDD B NET8 VDD P18 W=1.6U L=0.18U
MP4 NET8 D Z VDD P18 W=1.6U L=0.18U
MP2 NET8 E Z VDD P18 W=1.6U L=0.18U
MP1 VDD C NET8 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.6U L=0.18U
MN5 NET37 A GND GND N18 W=1.1U L=0.18U
MN6 NET45 D GND GND N18 W=1.0U L=0.18U
MN4 NET12 B NET37 GND N18 W=1.1U L=0.18U
MN1 Z C NET12 GND N18 W=1.1U L=0.18U
MN0 Z E NET45 GND N18 W=1.0U L=0.18U
.ENDS AOI32HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI31HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:31:17 2002                                       *
*******************************************************************************
.SUBCKT AOI31HDLX Z A B C D
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP2 NET8 D Z VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 Z C NET12 GND N18 W=0.58U L=0.18U
MN0 Z D GND GND N18 W=0.42U L=0.18U
.ENDS AOI31HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI31HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:31:16 2002                                       *
*******************************************************************************
.SUBCKT AOI31HD4X Z A B C D
XI4 NET27 NET54 IVG PW=1.6U NW=1.06U
XI5 Z NET27 IVG PW=4.8U NW=3.2U
MP3 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP2 NET8 D NET54 VDD P18 W=0.84U L=0.18U
MP1 VDD C NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN5 NET37 A GND GND N18 W=0.58U L=0.18U
MN4 NET12 B NET37 GND N18 W=0.58U L=0.18U
MN1 NET54 C NET12 GND N18 W=0.58U L=0.18U
MN0 NET54 D GND GND N18 W=0.42U L=0.18U
.ENDS AOI31HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI31HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:31:14 2002                                       *
*******************************************************************************
.SUBCKT AOI31HD2X Z A B C D
MP3 VDD B NET8 VDD P18 W=3.2U L=0.18U
MP2 NET8 D Z VDD P18 W=3.2U L=0.18U
MP1 VDD C NET8 VDD P18 W=3.2U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.2U L=0.18U
MN5 NET37 A GND GND N18 W=2.2U L=0.18U
MN4 NET12 B NET37 GND N18 W=2.2U L=0.18U
MN1 Z C NET12 GND N18 W=2.2U L=0.18U
MN0 Z D GND GND N18 W=1.6U L=0.18U
.ENDS AOI31HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI31HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:31:12 2002                                       *
*******************************************************************************
.SUBCKT AOI31HD1X Z A B C D
MP3 VDD B NET8 VDD P18 W=1.6U L=0.18U
MP2 NET8 D Z VDD P18 W=1.6U L=0.18U
MP1 VDD C NET8 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.6U L=0.18U
MN5 NET37 A GND GND N18 W=1.1U L=0.18U
MN4 NET12 B NET37 GND N18 W=1.1U L=0.18U
MN1 Z C NET12 GND N18 W=1.1U L=0.18U
MN0 Z D GND GND N18 W=0.8U L=0.18U
.ENDS AOI31HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:30:54 2002                                       *
*******************************************************************************
.SUBCKT AOI22HDLX Z A B C D
MP3 NET8 D Z VDD P18 W=0.84U L=0.18U
MP2 NET8 C Z VDD P18 W=0.84U L=0.18U
MP1 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN5 NET39 D GND GND N18 W=0.54U L=0.18U
MN4 NET12 A GND GND N18 W=0.54U L=0.18U
MN1 Z B NET12 GND N18 W=0.54U L=0.18U
MN0 Z C NET39 GND N18 W=0.54U L=0.18U
.ENDS AOI22HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:30:52 2002                                       *
*******************************************************************************
.SUBCKT AOI22HD4X Z A B C D
MP3 NET8 D Z VDD P18 W=6.4U L=0.18U
MP2 NET8 C Z VDD P18 W=6.4U L=0.18U
MP1 VDD B NET8 VDD P18 W=6.4U L=0.18U
MP0 VDD A NET8 VDD P18 W=6.4U L=0.18U
MN5 NET39 D GND GND N18 W=4.0U L=0.18U
MN4 NET12 A GND GND N18 W=4.0U L=0.18U
MN1 Z B NET12 GND N18 W=4.0U L=0.18U
MN0 Z C NET39 GND N18 W=4.0U L=0.18U
.ENDS AOI22HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:30:51 2002                                       *
*******************************************************************************
.SUBCKT AOI22HD2X Z A B C D
MP3 NET8 D Z VDD P18 W=3.2U L=0.18U
MP2 NET8 C Z VDD P18 W=3.2U L=0.18U
MP1 VDD B NET8 VDD P18 W=3.2U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.2U L=0.18U
MN5 NET39 D GND GND N18 W=2.0U L=0.18U
MN4 NET12 A GND GND N18 W=2.0U L=0.18U
MN1 Z B NET12 GND N18 W=2.0U L=0.18U
MN0 Z C NET39 GND N18 W=2.0U L=0.18U
.ENDS AOI22HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:30:49 2002                                       *
*******************************************************************************
.SUBCKT AOI22HD1X Z A B C D
MP3 NET8 D Z VDD P18 W=1.6U L=0.18U
MP2 NET8 C Z VDD P18 W=1.6U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.6U L=0.18U
MN5 NET39 D GND GND N18 W=1.0U L=0.18U
MN4 NET12 A GND GND N18 W=1.0U L=0.18U
MN1 Z B NET12 GND N18 W=1.0U L=0.18U
MN0 Z C NET39 GND N18 W=1.0U L=0.18U
.ENDS AOI22HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22B2HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:31:10 2002                                       *
*******************************************************************************
.SUBCKT AOI22B2HDLX Z AN BN C D
MP5 NET34 NET39 Z VDD P18 W=0.84U L=0.18U
MP4 VDD D NET34 VDD P18 W=0.84U L=0.18U
MP3 NET8 BN NET39 VDD P18 W=0.84U L=0.18U
MP2 VDD C NET34 VDD P18 W=0.84U L=0.18U
MP0 VDD AN NET8 VDD P18 W=0.84U L=0.18U
MN5 NET39 BN GND GND N18 W=0.42U L=0.18U
MN6 Z NET39 GND GND N18 W=0.42U L=0.18U
MN4 NET12 C GND GND N18 W=0.52U L=0.18U
MN1 Z D NET12 GND N18 W=0.52U L=0.18U
MN0 NET39 AN GND GND N18 W=0.42U L=0.18U
.ENDS AOI22B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22B2HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:31:08 2002                                       *
*******************************************************************************
.SUBCKT AOI22B2HD4X Z AN BN C D
MP5 NET34 NET39 Z VDD P18 W=6.4U L=0.18U
MP4 VDD D NET34 VDD P18 W=6.4U L=0.18U
MP3 NET8 BN NET39 VDD P18 W=1.68U L=0.18U
MP2 VDD C NET34 VDD P18 W=6.4U L=0.18U
MP0 VDD AN NET8 VDD P18 W=1.68U L=0.18U
MN5 NET39 BN GND GND N18 W=0.84U L=0.18U
MN6 Z NET39 GND GND N18 W=3.2U L=0.18U
MN4 NET12 C GND GND N18 W=4.0U L=0.18U
MN1 Z D NET12 GND N18 W=4.0U L=0.18U
MN0 NET39 AN GND GND N18 W=0.84U L=0.18U
.ENDS AOI22B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22B2HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:31:06 2002                                       *
*******************************************************************************
.SUBCKT AOI22B2HD2X Z AN BN C D
MP5 NET34 NET39 Z VDD P18 W=3.2U L=0.18U
MP4 VDD D NET34 VDD P18 W=3.2U L=0.18U
MP3 NET8 BN NET39 VDD P18 W=1.4U L=0.18U
MP2 VDD C NET34 VDD P18 W=3.2U L=0.18U
MP0 VDD AN NET8 VDD P18 W=1.4U L=0.18U
MN5 NET39 BN GND GND N18 W=0.7U L=0.18U
MN6 Z NET39 GND GND N18 W=1.6U L=0.18U
MN4 NET12 C GND GND N18 W=2.0U L=0.18U
MN1 Z D NET12 GND N18 W=2.0U L=0.18U
MN0 NET39 AN GND GND N18 W=0.7U L=0.18U
.ENDS AOI22B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI22B2HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:31:02 2002                                       *
*******************************************************************************
.SUBCKT AOI22B2HD1X Z AN BN C D
MP5 NET34 NET39 Z VDD P18 W=1.6U L=0.18U
MP4 VDD D NET34 VDD P18 W=1.6U L=0.18U
MP3 NET8 BN NET39 VDD P18 W=0.84U L=0.18U
MP2 VDD C NET34 VDD P18 W=1.6U L=0.18U
MP0 VDD AN NET8 VDD P18 W=0.84U L=0.18U
MN5 NET39 BN GND GND N18 W=0.42U L=0.18U
MN6 Z NET39 GND GND N18 W=0.8U L=0.18U
MN4 NET12 C GND GND N18 W=1.0U L=0.18U
MN1 Z D NET12 GND N18 W=1.0U L=0.18U
MN0 NET39 AN GND GND N18 W=0.42U L=0.18U
.ENDS AOI22B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI222HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:30:47 2002                                       *
*******************************************************************************
.SUBCKT AOI222HDLX Z A B C D E F
MP3 NET25 F Z VDD P18 W=0.98U L=0.18U
MP6 NET25 E Z VDD P18 W=0.98U L=0.18U
MP5 NET8 C NET25 VDD P18 W=0.98U L=0.18U
MP2 NET8 D NET25 VDD P18 W=0.98U L=0.18U
MP1 VDD B NET8 VDD P18 W=0.98U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.98U L=0.18U
MN7 NET55 E GND GND N18 W=0.52U L=0.18U
MN6 NET43 C GND GND N18 W=0.52U L=0.18U
MN5 Z D NET43 GND N18 W=0.52U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 Z B NET12 GND N18 W=0.52U L=0.18U
MN0 Z F NET55 GND N18 W=0.52U L=0.18U
.ENDS AOI222HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI222HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:30:46 2002                                       *
*******************************************************************************
.SUBCKT AOI222HD4X Z A B C D E F
XI4 NET40 NET76 IVG PW=1.6U NW=1.06U
XI5 Z NET40 IVG PW=4.8U NW=3.2U
MP3 NET25 F NET76 VDD P18 W=1.0U L=0.18U
MP6 NET25 E NET76 VDD P18 W=1.0U L=0.18U
MP5 NET8 C NET25 VDD P18 W=1.0U L=0.18U
MP2 NET8 D NET25 VDD P18 W=1.0U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.0U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.0U L=0.18U
MN7 NET55 E GND GND N18 W=0.52U L=0.18U
MN6 NET43 C GND GND N18 W=0.52U L=0.18U
MN5 NET76 D NET43 GND N18 W=0.52U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 NET76 B NET12 GND N18 W=0.52U L=0.18U
MN0 NET76 F NET55 GND N18 W=0.52U L=0.18U
.ENDS AOI222HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI222HD2X                                                           *
* LAST TIME SAVED: JUL 14 11:20:36 2004                                       *
*******************************************************************************
.SUBCKT AOI222HD2X Z A B C D E F
XI4 NET40 NET76 IVG PW=0.8U NW=0.53U
XI5 Z NET40 IVG PW=2.4U NW=1.6U
MP3 NET25 F NET76 VDD P18 W=0.81U L=0.18U
MP6 NET25 E NET76 VDD P18 W=0.81U L=0.18U
MP5 NET8 C NET25 VDD P18 W=0.81U L=0.18U
MP2 NET8 D NET25 VDD P18 W=0.81U L=0.18U
MP1 VDD B NET8 VDD P18 W=0.81U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.81U L=0.18U
MN7 NET55 E GND GND N18 W=0.42U L=0.18U
MN6 NET43 C GND GND N18 W=0.42U L=0.18U
MN5 NET76 D NET43 GND N18 W=0.42U L=0.18U
MN4 NET12 A GND GND N18 W=0.42U L=0.18U
MN1 NET76 B NET12 GND N18 W=0.42U L=0.18U
MN0 NET76 F NET55 GND N18 W=0.42U L=0.18U
.ENDS AOI222HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI222HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:30:42 2002                                       *
*******************************************************************************
.SUBCKT AOI222HD1X Z A B C D E F
MP3 NET25 F Z VDD P18 W=1.68U L=0.18U
MP6 NET25 E Z VDD P18 W=1.68U L=0.18U
MP5 NET8 C NET25 VDD P18 W=1.68U L=0.18U
MP2 NET8 D NET25 VDD P18 W=1.68U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.68U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.68U L=0.18U
MN7 NET55 E GND GND N18 W=0.88U L=0.18U
MN6 NET43 C GND GND N18 W=0.88U L=0.18U
MN5 Z D NET43 GND N18 W=0.88U L=0.18U
MN4 NET12 A GND GND N18 W=0.88U L=0.18U
MN1 Z B NET12 GND N18 W=0.88U L=0.18U
MN0 Z F NET55 GND N18 W=0.88U L=0.18U
.ENDS AOI222HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI221HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:30:40 2002                                       *
*******************************************************************************
.SUBCKT AOI221HDLX Z A B C D E
MP3 NET25 E Z VDD P18 W=1.0U L=0.18U
MP5 NET8 C NET25 VDD P18 W=1.0U L=0.18U
MP2 NET8 D NET25 VDD P18 W=1.0U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.0U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.0U L=0.18U
MN6 NET43 C GND GND N18 W=0.52U L=0.18U
MN5 Z D NET43 GND N18 W=0.52U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 Z B NET12 GND N18 W=0.52U L=0.18U
MN0 Z E GND GND N18 W=0.42U L=0.18U
.ENDS AOI221HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI221HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:30:38 2002                                       *
*******************************************************************************
.SUBCKT AOI221HD4X Z A B C D E
XI4 NET34 NET64 IVG PW=1.6U NW=1.06U
XI5 Z NET34 IVG PW=4.8U NW=3.2U
MP3 NET25 E NET64 VDD P18 W=1.0U L=0.18U
MP5 NET8 C NET25 VDD P18 W=1.0U L=0.18U
MP2 NET8 D NET25 VDD P18 W=1.0U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.0U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.0U L=0.18U
MN6 NET43 C GND GND N18 W=0.52U L=0.18U
MN5 NET64 D NET43 GND N18 W=0.52U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 NET64 B NET12 GND N18 W=0.52U L=0.18U
MN0 NET64 E GND GND N18 W=0.42U L=0.18U
.ENDS AOI221HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI221HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:30:37 2002                                       *
*******************************************************************************
.SUBCKT AOI221HD2X Z A B C D E
MP3 NET25 E Z VDD P18 W=3.36U L=0.18U
MP5 NET8 C NET25 VDD P18 W=3.36U L=0.18U
MP2 NET8 D NET25 VDD P18 W=3.36U L=0.18U
MP1 VDD B NET8 VDD P18 W=3.36U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.36U L=0.18U
MN6 NET43 C GND GND N18 W=1.76U L=0.18U
MN5 Z D NET43 GND N18 W=1.76U L=0.18U
MN4 NET12 A GND GND N18 W=1.76U L=0.18U
MN1 Z B NET12 GND N18 W=1.76U L=0.18U
MN0 Z E GND GND N18 W=1.4U L=0.18U
.ENDS AOI221HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI221HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:30:35 2002                                       *
*******************************************************************************
.SUBCKT AOI221HD1X Z A B C D E
MP3 NET25 E Z VDD P18 W=1.68U L=0.18U
MP5 NET8 C NET25 VDD P18 W=1.68U L=0.18U
MP2 NET8 D NET25 VDD P18 W=1.68U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.68U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.68U L=0.18U
MN6 NET43 C GND GND N18 W=0.88U L=0.18U
MN5 Z D NET43 GND N18 W=0.88U L=0.18U
MN4 NET12 A GND GND N18 W=0.88U L=0.18U
MN1 Z B NET12 GND N18 W=0.88U L=0.18U
MN0 Z E GND GND N18 W=0.7U L=0.18U
.ENDS AOI221HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21HDLX                                                            *
* LAST TIME SAVED: AUG 30 10:30:34 2002                                       *
*******************************************************************************
.SUBCKT AOI21HDLX Z A B C
MP2 NET8 C Z VDD P18 W=0.84U L=0.18U
MP1 VDD B NET8 VDD P18 W=0.84U L=0.18U
MP0 VDD A NET8 VDD P18 W=0.84U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 Z B NET12 GND N18 W=0.52U L=0.18U
MN0 Z C GND GND N18 W=0.42U L=0.18U
.ENDS AOI21HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21HD4X                                                            *
* LAST TIME SAVED: AUG 30 10:30:32 2002                                       *
*******************************************************************************
.SUBCKT AOI21HD4X Z A B C
MP2 NET8 C Z VDD P18 W=6.4U L=0.18U
MP1 VDD B NET8 VDD P18 W=6.4U L=0.18U
MP0 VDD A NET8 VDD P18 W=6.4U L=0.18U
MN4 NET12 A GND GND N18 W=4.0U L=0.18U
MN1 Z B NET12 GND N18 W=4.0U L=0.18U
MN0 Z C GND GND N18 W=3.2U L=0.18U
.ENDS AOI21HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21HD2X                                                            *
* LAST TIME SAVED: AUG 30 10:30:30 2002                                       *
*******************************************************************************
.SUBCKT AOI21HD2X Z A B C
MP2 NET8 C Z VDD P18 W=3.2U L=0.18U
MP1 VDD B NET8 VDD P18 W=3.2U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.2U L=0.18U
MN4 NET12 A GND GND N18 W=2.0U L=0.18U
MN1 Z B NET12 GND N18 W=2.0U L=0.18U
MN0 Z C GND GND N18 W=1.6U L=0.18U
.ENDS AOI21HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21HD1X                                                            *
* LAST TIME SAVED: AUG 30 10:30:28 2002                                       *
*******************************************************************************
.SUBCKT AOI21HD1X Z A B C
MP2 NET8 C Z VDD P18 W=1.6U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.6U L=0.18U
MN4 NET12 A GND GND N18 W=1.0U L=0.18U
MN1 Z B NET12 GND N18 W=1.0U L=0.18U
MN0 Z C GND GND N18 W=0.8U L=0.18U
.ENDS AOI21HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21B2HDLX                                                          *
* LAST TIME SAVED: AUG 30 10:31:00 2002                                       *
*******************************************************************************
.SUBCKT AOI21B2HDLX Z AN BN C
MP3 VDD AN NET28 VDD P18 W=0.84U L=0.18U
MP4 NET28 BN NET22 VDD P18 W=0.84U L=0.18U
MP2 NET8 C Z VDD P18 W=0.84U L=0.18U
MP1 VDD NET22 NET8 VDD P18 W=0.84U L=0.18U
MN5 NET22 AN GND GND N18 W=0.42U L=0.18U
MN4 Z C GND GND N18 W=0.42U L=0.18U
MN7 Z NET22 GND GND N18 W=0.42U L=0.18U
MN6 NET22 BN GND GND N18 W=0.42U L=0.18U
.ENDS AOI21B2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21B2HD4X                                                          *
* LAST TIME SAVED: AUG 30 10:30:59 2002                                       *
*******************************************************************************
.SUBCKT AOI21B2HD4X Z AN BN C
MP3 VDD AN NET28 VDD P18 W=1.68U L=0.18U
MP4 NET28 BN NET22 VDD P18 W=1.68U L=0.18U
MP2 NET8 C Z VDD P18 W=6.4U L=0.18U
MP1 VDD NET22 NET8 VDD P18 W=6.4U L=0.18U
MN5 NET22 AN GND GND N18 W=0.84U L=0.18U
MN4 Z C GND GND N18 W=3.2U L=0.18U
MN7 Z NET22 GND GND N18 W=3.2U L=0.18U
MN6 NET22 BN GND GND N18 W=0.84U L=0.18U
.ENDS AOI21B2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21B2HD2X                                                          *
* LAST TIME SAVED: AUG 30 10:30:57 2002                                       *
*******************************************************************************
.SUBCKT AOI21B2HD2X Z AN BN C
MP3 VDD AN NET28 VDD P18 W=1.4U L=0.18U
MP4 NET28 BN NET22 VDD P18 W=1.4U L=0.18U
MP2 NET8 C Z VDD P18 W=3.2U L=0.18U
MP1 VDD NET22 NET8 VDD P18 W=3.2U L=0.18U
MN5 NET22 AN GND GND N18 W=0.7U L=0.18U
MN4 Z C GND GND N18 W=1.6U L=0.18U
MN7 Z NET22 GND GND N18 W=1.6U L=0.18U
MN6 NET22 BN GND GND N18 W=0.7U L=0.18U
.ENDS AOI21B2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI21B2HD1X                                                          *
* LAST TIME SAVED: AUG 30 10:30:55 2002                                       *
*******************************************************************************
.SUBCKT AOI21B2HD1X Z AN BN C
MP3 VDD AN NET28 VDD P18 W=0.84U L=0.18U
MP4 NET28 BN NET22 VDD P18 W=0.84U L=0.18U
MP2 NET8 C Z VDD P18 W=1.6U L=0.18U
MP1 VDD NET22 NET8 VDD P18 W=1.6U L=0.18U
MN5 NET22 AN GND GND N18 W=0.42U L=0.18U
MN4 Z C GND GND N18 W=0.8U L=0.18U
MN7 Z NET22 GND GND N18 W=0.8U L=0.18U
MN6 NET22 BN GND GND N18 W=0.42U L=0.18U
.ENDS AOI21B2HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI211HDLX                                                           *
* LAST TIME SAVED: AUG 30 10:30:26 2002                                       *
*******************************************************************************
.SUBCKT AOI211HDLX Z A B C D
MP3 NET25 D Z VDD P18 W=1.0U L=0.18U
MP2 NET8 C NET25 VDD P18 W=1.0U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.0U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.0U L=0.18U
MN5 Z D GND GND N18 W=0.42U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 Z B NET12 GND N18 W=0.52U L=0.18U
MN0 Z C GND GND N18 W=0.42U L=0.18U
.ENDS AOI211HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI211HD4X                                                           *
* LAST TIME SAVED: AUG 30 10:30:24 2002                                       *
*******************************************************************************
.SUBCKT AOI211HD4X Z A B C D
XI4 NET54 NET52 IVG PW=1.6U NW=1.06U
XI5 Z NET54 IVG PW=4.8U NW=3.2U
MP3 NET25 D NET52 VDD P18 W=1.0U L=0.18U
MP2 NET8 C NET25 VDD P18 W=1.0U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.0U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.0U L=0.18U
MN5 NET52 D GND GND N18 W=0.42U L=0.18U
MN4 NET12 A GND GND N18 W=0.52U L=0.18U
MN1 NET52 B NET12 GND N18 W=0.52U L=0.18U
MN0 NET52 C GND GND N18 W=0.42U L=0.18U
.ENDS AOI211HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI211HD2X                                                           *
* LAST TIME SAVED: AUG 30 10:30:22 2002                                       *
*******************************************************************************
.SUBCKT AOI211HD2X Z A B C D
MP3 NET25 D Z VDD P18 W=3.36U L=0.18U
MP2 NET8 C NET25 VDD P18 W=3.36U L=0.18U
MP1 VDD B NET8 VDD P18 W=3.36U L=0.18U
MP0 VDD A NET8 VDD P18 W=3.36U L=0.18U
MN5 Z D GND GND N18 W=1.4U L=0.18U
MN4 NET12 A GND GND N18 W=1.76U L=0.18U
MN1 Z B NET12 GND N18 W=1.76U L=0.18U
MN0 Z C GND GND N18 W=1.4U L=0.18U
.ENDS AOI211HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AOI211HD1X                                                           *
* LAST TIME SAVED: AUG 30 10:30:20 2002                                       *
*******************************************************************************
.SUBCKT AOI211HD1X Z A B C D
MP3 NET25 D Z VDD P18 W=1.68U L=0.18U
MP2 NET8 C NET25 VDD P18 W=1.68U L=0.18U
MP1 VDD B NET8 VDD P18 W=1.68U L=0.18U
MP0 VDD A NET8 VDD P18 W=1.68U L=0.18U
MN5 Z D GND GND N18 W=0.7U L=0.18U
MN4 NET12 A GND GND N18 W=0.88U L=0.18U
MN1 Z B NET12 GND N18 W=0.88U L=0.18U
MN0 Z C GND GND N18 W=0.7U L=0.18U
.ENDS AOI211HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: ANTFIXHD                                                             *
* LAST TIME SAVED: DEC 16 10:36:40 2003                                       *
*******************************************************************************
.SUBCKT ANTFIXHD Z
*.NOPIN VDD
D0 GND Z NDIO18 AREA=1.086P W=1.04U L=1.04U
.ENDS ANTFIXHD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND4HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:30:18 2002                                       *
*******************************************************************************
.SUBCKT AND4HDLX Z A B C D
XI3 Z NET35 IVG PW=0.64U NW=0.42U
MN4 NET7 B NET28 GND N18 W=0.64U L=0.18U
MN5 NET28 A GND GND N18 W=0.64U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.64U L=0.18U
MN0 NET35 D NET10 GND N18 W=0.64U L=0.18U
MP3 VDD A NET35 VDD P18 W=0.64U L=0.18U
MP2 VDD D NET35 VDD P18 W=0.64U L=0.18U
MP1 VDD C NET35 VDD P18 W=0.64U L=0.18U
MP0 VDD B NET35 VDD P18 W=0.64U L=0.18U
.ENDS AND4HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND4HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:30:16 2002                                       *
*******************************************************************************
.SUBCKT AND4HD4X Z A B C D
XI3 Z NET35 IVG PW=4.8U NW=3.2U
MN4 NET7 B NET28 GND N18 W=1.18U L=0.18U
MN5 NET28 A GND GND N18 W=1.18U L=0.18U
MN3 NET10 C NET7 GND N18 W=1.18U L=0.18U
MN0 NET35 D NET10 GND N18 W=1.18U L=0.18U
MP3 VDD A NET35 VDD P18 W=1.18U L=0.18U
MP2 VDD D NET35 VDD P18 W=1.18U L=0.18U
MP1 VDD C NET35 VDD P18 W=1.18U L=0.18U
MP0 VDD B NET35 VDD P18 W=1.18U L=0.18U
.ENDS AND4HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND4HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:30:14 2002                                       *
*******************************************************************************
.SUBCKT AND4HD2X Z A B C D
XI3 Z NET35 IVG PW=2.4U NW=1.6U
MN4 NET7 B NET28 GND N18 W=0.8U L=0.18U
MN5 NET28 A GND GND N18 W=0.8U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.8U L=0.18U
MN0 NET35 D NET10 GND N18 W=0.8U L=0.18U
MP3 VDD A NET35 VDD P18 W=0.8U L=0.18U
MP2 VDD D NET35 VDD P18 W=0.8U L=0.18U
MP1 VDD C NET35 VDD P18 W=0.8U L=0.18U
MP0 VDD B NET35 VDD P18 W=0.8U L=0.18U
.ENDS AND4HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND4HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:30:12 2002                                       *
*******************************************************************************
.SUBCKT AND4HD1X Z A B C D
XI3 Z NET35 IVG PW=1.2U NW=0.8U
MN4 NET7 B NET59 GND N18 W=0.64U L=0.18U
MN5 NET59 A GND GND N18 W=0.64U L=0.18U
MN3 NET10 C NET7 GND N18 W=0.64U L=0.18U
MN0 NET35 D NET10 GND N18 W=0.64U L=0.18U
MP3 VDD A NET35 VDD P18 W=0.64U L=0.18U
MP2 VDD D NET35 VDD P18 W=0.64U L=0.18U
MP1 VDD C NET35 VDD P18 W=0.64U L=0.18U
MP0 VDD B NET35 VDD P18 W=0.64U L=0.18U
.ENDS AND4HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND3HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:30:10 2002                                       *
*******************************************************************************
.SUBCKT AND3HDLX Z A B C
XI2 Z NET36 IVG PW=0.64U NW=0.42U
MN4 NET7 A GND GND N18 W=0.58U L=0.18U
MN3 NET10 B NET7 GND N18 W=0.58U L=0.18U
MN0 NET36 C NET10 GND N18 W=0.58U L=0.18U
MP2 VDD C NET36 VDD P18 W=0.64U L=0.18U
MP1 VDD B NET36 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET36 VDD P18 W=0.64U L=0.18U
.ENDS AND3HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND3HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:30:08 2002                                       *
*******************************************************************************
.SUBCKT AND3HD4X Z A B C
XI2 Z NET36 IVG PW=4.8U NW=3.2U
MN4 NET7 A GND GND N18 W=1.18U L=0.18U
MN3 NET10 B NET7 GND N18 W=1.18U L=0.18U
MN0 NET36 C NET10 GND N18 W=1.18U L=0.18U
MP2 VDD C NET36 VDD P18 W=1.6U L=0.18U
MP1 VDD B NET36 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET36 VDD P18 W=1.6U L=0.18U
.ENDS AND3HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND3HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:30:07 2002                                       *
*******************************************************************************
.SUBCKT AND3HD2X Z A B C
XI2 Z NET36 IVG PW=2.4U NW=1.6U
MN4 NET7 A GND GND N18 W=0.74U L=0.18U
MN3 NET10 B NET7 GND N18 W=0.74U L=0.18U
MN0 NET36 C NET10 GND N18 W=0.74U L=0.18U
MP2 VDD C NET36 VDD P18 W=0.8U L=0.18U
MP1 VDD B NET36 VDD P18 W=0.8U L=0.18U
MP0 VDD A NET36 VDD P18 W=0.8U L=0.18U
.ENDS AND3HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND3HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:30:06 2002                                       *
*******************************************************************************
.SUBCKT AND3HD1X Z A B C
XI2 Z NET36 IVG PW=1.2U NW=0.8U
MN4 NET7 A GND GND N18 W=0.58U L=0.18U
MN3 NET10 B NET7 GND N18 W=0.58U L=0.18U
MN0 NET36 C NET10 GND N18 W=0.58U L=0.18U
MP2 VDD C NET36 VDD P18 W=0.64U L=0.18U
MP1 VDD B NET36 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET36 VDD P18 W=0.64U L=0.18U
.ENDS AND3HD1X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HDLX                                                             *
* LAST TIME SAVED: AUG 30 10:30:03 2002                                       *
*******************************************************************************
.SUBCKT AND2HDLX Z A B
XI2 Z NET26 IVG PW=0.64U NW=0.42U
MN1 NET6 A GND GND N18 W=0.54U L=0.18U
MN0 NET26 B NET6 GND N18 W=0.54U L=0.18U
MP1 VDD B NET26 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET26 VDD P18 W=0.64U L=0.18U
.ENDS AND2HDLX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HD4XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:30:02 2002                                       *
*******************************************************************************
.SUBCKT AND2HD4XSPG Z A B
XI2 Z NET26 IVG PW=4.8U NW=3.2U
MN1 NET6 A GND GND N18 W=1.18U L=0.18U
MN0 NET26 B NET6 GND N18 W=1.18U L=0.18U
MP1 VDD B NET26 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET26 VDD P18 W=1.6U L=0.18U
.ENDS AND2HD4XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HD4X                                                             *
* LAST TIME SAVED: AUG 30 10:30:01 2002                                       *
*******************************************************************************
.SUBCKT AND2HD4X Z A B
XI2 Z NET26 IVG PW=4.8U NW=3.2U
MN1 NET6 A GND GND N18 W=1.18U L=0.18U
MN0 NET26 B NET6 GND N18 W=1.18U L=0.18U
MP1 VDD B NET26 VDD P18 W=1.6U L=0.18U
MP0 VDD A NET26 VDD P18 W=1.6U L=0.18U
.ENDS AND2HD4X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HD2XSPG                                                          *
* LAST TIME SAVED: AUG 30 10:30:00 2002                                       *
*******************************************************************************
.SUBCKT AND2HD2XSPG Z A B
XI2 Z NET26 IVG PW=2.4U NW=1.6U
MN1 NET6 A GND GND N18 W=0.66U L=0.18U
MN0 NET26 B NET6 GND N18 W=0.66U L=0.18U
MP1 VDD B NET26 VDD P18 W=0.8U L=0.18U
MP0 VDD A NET26 VDD P18 W=0.8U L=0.18U
.ENDS AND2HD2XSPG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HD2X                                                             *
* LAST TIME SAVED: AUG 30 10:29:53 2002                                       *
*******************************************************************************
.SUBCKT AND2HD2X Z A B
XI2 Z NET26 IVG PW=2.4U NW=1.6U
MN1 NET6 A GND GND N18 W=0.66U L=0.18U
MN0 NET26 B NET6 GND N18 W=0.66U L=0.18U
MP1 VDD B NET26 VDD P18 W=0.8U L=0.18U
MP0 VDD A NET26 VDD P18 W=0.8U L=0.18U
.ENDS AND2HD2X


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AND2HD1X                                                             *
* LAST TIME SAVED: AUG 30 10:29:51 2002                                       *
*******************************************************************************
.SUBCKT AND2HD1X Z A B
XI2 Z NET26 IVG PW=1.2U NW=0.8U
MN1 NET6 A GND GND N18 W=0.54U L=0.18U
MN0 NET26 B NET6 GND N18 W=0.54U L=0.18U
MP1 VDD B NET26 VDD P18 W=0.64U L=0.18U
MP0 VDD A NET26 VDD P18 W=0.64U L=0.18U
.ENDS AND2HD1X
